module PositPackedtoUnpacked(
  input         clock,
  input         reset,
  input         io_in_sign,
  input  [14:0] io_in_others,
  output        io_out_sign,
  output [27:0] io_out_exponent,
  output [11:0] io_out_fraction
);
  wire [14:0] _T_1; // @[Bitwise.scala 71:12]
  wire [14:0] _T_2; // @[Conversion.scala 15:36]
  wire [14:0] _GEN_0; // @[Conversion.scala 15:79]
  wire [14:0] others; // @[Conversion.scala 15:79]
  wire [14:0] _T_5; // @[Conversion.scala 16:129]
  wire [7:0] _T_10; // @[Bitwise.scala 102:31]
  wire [7:0] _T_12; // @[Bitwise.scala 102:65]
  wire [7:0] _T_14; // @[Bitwise.scala 102:75]
  wire [7:0] _T_15; // @[Bitwise.scala 102:39]
  wire [7:0] _GEN_1; // @[Bitwise.scala 102:31]
  wire [7:0] _T_20; // @[Bitwise.scala 102:31]
  wire [7:0] _T_22; // @[Bitwise.scala 102:65]
  wire [7:0] _T_24; // @[Bitwise.scala 102:75]
  wire [7:0] _T_25; // @[Bitwise.scala 102:39]
  wire [7:0] _GEN_2; // @[Bitwise.scala 102:31]
  wire [7:0] _T_30; // @[Bitwise.scala 102:31]
  wire [7:0] _T_32; // @[Bitwise.scala 102:65]
  wire [7:0] _T_34; // @[Bitwise.scala 102:75]
  wire [7:0] _T_35; // @[Bitwise.scala 102:39]
  wire [14:0] _T_55; // @[Cat.scala 29:58]
  wire [3:0] _T_71; // @[Mux.scala 47:69]
  wire [3:0] _T_72; // @[Mux.scala 47:69]
  wire [3:0] _T_73; // @[Mux.scala 47:69]
  wire [3:0] _T_74; // @[Mux.scala 47:69]
  wire [3:0] _T_75; // @[Mux.scala 47:69]
  wire [3:0] _T_76; // @[Mux.scala 47:69]
  wire [3:0] _T_77; // @[Mux.scala 47:69]
  wire [3:0] _T_78; // @[Mux.scala 47:69]
  wire [3:0] _T_79; // @[Mux.scala 47:69]
  wire [3:0] _T_80; // @[Mux.scala 47:69]
  wire [3:0] _T_81; // @[Mux.scala 47:69]
  wire [3:0] _T_82; // @[Mux.scala 47:69]
  wire [3:0] _T_83; // @[Mux.scala 47:69]
  wire [3:0] leading; // @[Mux.scala 47:69]
  assign _T_1 = io_in_sign ? 15'h7fff : 15'h0; // @[Bitwise.scala 71:12]
  assign _T_2 = io_in_others ^ _T_1; // @[Conversion.scala 15:36]
  assign _GEN_0 = {{14'd0}, io_in_sign}; // @[Conversion.scala 15:79]
  assign others = _T_2 + _GEN_0; // @[Conversion.scala 15:79]
  assign _T_5 = ~others; // @[Conversion.scala 16:129]
  assign _T_10 = {{4'd0}, _T_5[7:4]}; // @[Bitwise.scala 102:31]
  assign _T_12 = {_T_5[3:0], 4'h0}; // @[Bitwise.scala 102:65]
  assign _T_14 = _T_12 & 8'hf0; // @[Bitwise.scala 102:75]
  assign _T_15 = _T_10 | _T_14; // @[Bitwise.scala 102:39]
  assign _GEN_1 = {{2'd0}, _T_15[7:2]}; // @[Bitwise.scala 102:31]
  assign _T_20 = _GEN_1 & 8'h33; // @[Bitwise.scala 102:31]
  assign _T_22 = {_T_15[5:0], 2'h0}; // @[Bitwise.scala 102:65]
  assign _T_24 = _T_22 & 8'hcc; // @[Bitwise.scala 102:75]
  assign _T_25 = _T_20 | _T_24; // @[Bitwise.scala 102:39]
  assign _GEN_2 = {{1'd0}, _T_25[7:1]}; // @[Bitwise.scala 102:31]
  assign _T_30 = _GEN_2 & 8'h55; // @[Bitwise.scala 102:31]
  assign _T_32 = {_T_25[6:0], 1'h0}; // @[Bitwise.scala 102:65]
  assign _T_34 = _T_32 & 8'haa; // @[Bitwise.scala 102:75]
  assign _T_35 = _T_30 | _T_34; // @[Bitwise.scala 102:39]
  assign _T_55 = {_T_35,_T_5[8],_T_5[9],_T_5[10],_T_5[11],_T_5[12],_T_5[13],_T_5[14]}; // @[Cat.scala 29:58]
  assign _T_71 = _T_55[13] ? 4'hd : 4'he; // @[Mux.scala 47:69]
  assign _T_72 = _T_55[12] ? 4'hc : _T_71; // @[Mux.scala 47:69]
  assign _T_73 = _T_55[11] ? 4'hb : _T_72; // @[Mux.scala 47:69]
  assign _T_74 = _T_55[10] ? 4'ha : _T_73; // @[Mux.scala 47:69]
  assign _T_75 = _T_55[9] ? 4'h9 : _T_74; // @[Mux.scala 47:69]
  assign _T_76 = _T_55[8] ? 4'h8 : _T_75; // @[Mux.scala 47:69]
  assign _T_77 = _T_55[7] ? 4'h7 : _T_76; // @[Mux.scala 47:69]
  assign _T_78 = _T_55[6] ? 4'h6 : _T_77; // @[Mux.scala 47:69]
  assign _T_79 = _T_55[5] ? 4'h5 : _T_78; // @[Mux.scala 47:69]
  assign _T_80 = _T_55[4] ? 4'h4 : _T_79; // @[Mux.scala 47:69]
  assign _T_81 = _T_55[3] ? 4'h3 : _T_80; // @[Mux.scala 47:69]
  assign _T_82 = _T_55[2] ? 4'h2 : _T_81; // @[Mux.scala 47:69]
  assign _T_83 = _T_55[1] ? 4'h1 : _T_82; // @[Mux.scala 47:69]
  assign leading = _T_55[0] ? 4'h0 : _T_83; // @[Mux.scala 47:69]
  assign io_out_sign = io_in_sign; // @[Conversion.scala 13:21]
  assign io_out_exponent = {{24'd0}, leading}; // @[Conversion.scala 17:25]
  assign io_out_fraction = 12'h0; // @[Conversion.scala 18:25]
endmodule
