module logMultiplier(
  input          io_A_zero,
  input          io_A_nan,
  input          io_A_sign,
  input  [5:0]   io_A_exponent,
  input  [12:0]  io_A_fraction,
  input          io_B_zero,
  input          io_B_nan,
  input          io_B_sign,
  input  [5:0]   io_B_exponent,
  input  [12:0]  io_B_fraction,
  output         io_out_zero,
  output         io_out_nan,
  output [128:0] io_out_number
);
  wire [6:0] exponentSum; // @[Multiplier.scala 60:49]
  wire [12:0] fractionSum; // @[Multiplier.scala 61:71]
  wire [7:0] _T_4; // @[Multiplier.scala 63:42]
  wire [8:0] shift; // @[Multiplier.scala 63:57]
  wire  _T_5; // @[Multiplier.scala 64:32]
  wire [8:0] _T_9; // @[Multiplier.scala 64:67]
  wire [9:0] _GEN_3; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_4; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_5; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_6; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_7; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_8; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_9; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_10; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_11; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_12; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_13; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_14; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_15; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_16; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_17; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_18; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_19; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_20; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_21; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_22; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_23; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_24; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_25; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_26; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_27; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_28; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_29; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_30; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_31; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_32; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_33; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_34; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_35; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_36; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_37; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_38; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_39; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_40; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_41; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_42; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_43; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_44; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_45; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_46; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_47; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_48; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_49; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_50; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_51; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_52; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_53; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_54; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_55; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_56; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_57; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_58; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_59; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_60; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_61; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_62; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_63; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_64; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_65; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_66; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_67; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_68; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_69; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_70; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_71; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_72; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_73; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_74; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_75; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_76; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_77; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_78; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_79; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_80; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_81; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_82; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_83; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_84; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_85; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_86; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_87; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_88; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_89; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_90; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_91; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_92; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_93; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_94; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_95; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_96; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_97; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_98; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_99; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_100; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_101; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_102; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_103; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_104; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_105; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_106; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_107; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_108; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_109; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_110; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_111; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_112; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_113; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_114; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_115; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_116; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_117; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_118; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_119; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_120; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_121; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_122; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_123; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_124; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_125; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_126; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_127; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_128; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_129; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_130; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_131; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_132; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_133; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_134; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_135; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_136; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_137; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_138; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_139; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_140; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_141; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_142; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_143; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_144; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_145; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_146; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_147; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_148; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_149; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_150; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_151; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_152; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_153; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_154; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_155; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_156; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_157; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_158; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_159; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_160; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_161; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_162; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_163; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_164; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_165; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_166; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_167; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_168; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_169; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_170; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_171; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_172; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_173; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_174; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_175; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_176; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_177; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_178; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_179; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_180; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_181; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_182; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_183; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_184; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_185; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_186; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_187; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_188; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_189; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_190; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_191; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_192; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_193; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_194; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_195; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_196; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_197; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_198; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_199; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_200; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_201; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_202; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_203; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_204; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_205; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_206; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_207; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_208; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_209; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_210; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_211; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_212; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_213; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_214; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_215; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_216; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_217; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_218; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_219; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_220; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_221; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_222; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_223; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_224; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_225; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_226; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_227; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_228; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_229; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_230; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_231; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_232; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_233; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_234; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_235; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_236; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_237; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_238; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_239; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_240; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_241; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_242; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_243; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_244; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_245; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_246; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_247; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_248; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_249; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_250; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_251; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_252; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_253; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_254; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_255; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_256; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_257; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_258; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_259; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_260; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_261; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_262; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_263; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_264; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_265; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_266; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_267; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_268; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_269; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_270; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_271; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_272; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_273; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_274; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_275; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_276; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_277; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_278; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_279; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_280; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_281; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_282; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_283; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_284; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_285; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_286; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_287; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_288; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_289; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_290; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_291; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_292; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_293; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_294; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_295; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_296; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_297; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_298; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_299; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_300; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_301; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_302; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_303; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_304; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_305; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_306; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_307; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_308; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_309; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_310; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_311; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_312; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_313; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_314; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_315; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_316; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_317; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_318; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_319; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_320; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_321; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_322; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_323; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_324; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_325; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_326; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_327; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_328; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_329; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_330; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_331; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_332; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_333; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_334; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_335; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_336; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_337; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_338; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_339; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_340; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_341; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_342; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_343; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_344; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_345; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_346; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_347; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_348; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_349; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_350; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_351; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_352; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_353; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_354; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_355; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_356; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_357; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_358; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_359; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_360; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_361; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_362; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_363; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_364; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_365; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_366; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_367; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_368; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_369; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_370; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_371; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_372; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_373; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_374; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_375; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_376; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_377; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_378; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_379; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_380; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_381; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_382; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_383; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_384; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_385; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_386; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_387; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_388; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_389; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_390; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_391; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_392; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_393; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_394; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_395; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_396; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_397; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_398; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_399; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_400; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_401; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_402; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_403; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_404; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_405; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_406; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_407; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_408; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_409; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_410; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_411; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_412; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_413; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_414; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_415; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_416; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_417; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_418; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_419; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_420; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_421; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_422; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_423; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_424; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_425; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_426; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_427; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_428; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_429; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_430; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_431; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_432; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_433; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_434; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_435; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_436; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_437; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_438; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_439; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_440; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_441; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_442; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_443; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_444; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_445; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_446; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_447; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_448; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_449; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_450; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_451; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_452; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_453; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_454; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_455; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_456; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_457; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_458; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_459; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_460; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_461; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_462; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_463; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_464; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_465; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_466; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_467; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_468; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_469; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_470; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_471; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_472; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_473; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_474; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_475; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_476; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_477; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_478; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_479; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_480; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_481; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_482; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_483; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_484; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_485; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_486; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_487; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_488; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_489; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_490; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_491; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_492; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_493; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_494; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_495; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_496; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_497; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_498; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_499; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_500; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_501; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_502; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_503; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_504; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_505; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_506; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_507; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_508; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_509; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_510; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_511; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_512; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_513; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_514; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_515; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_516; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_517; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_518; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_519; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_520; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_521; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_522; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_523; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_524; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_525; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_526; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_527; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_528; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_529; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_530; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_531; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_532; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_533; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_534; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_535; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_536; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_537; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_538; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_539; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_540; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_541; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_542; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_543; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_544; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_545; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_546; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_547; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_548; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_549; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_550; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_551; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_552; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_553; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_554; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_555; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_556; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_557; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_558; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_559; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_560; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_561; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_562; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_563; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_564; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_565; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_566; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_567; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_568; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_569; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_570; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_571; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_572; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_573; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_574; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_575; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_576; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_577; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_578; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_579; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_580; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_581; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_582; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_583; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_584; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_585; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_586; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_587; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_588; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_589; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_590; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_591; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_592; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_593; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_594; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_595; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_596; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_597; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_598; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_599; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_600; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_601; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_602; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_603; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_604; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_605; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_606; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_607; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_608; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_609; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_610; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_611; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_612; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_613; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_614; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_615; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_616; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_617; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_618; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_619; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_620; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_621; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_622; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_623; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_624; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_625; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_626; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_627; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_628; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_629; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_630; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_631; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_632; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_633; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_634; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_635; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_636; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_637; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_638; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_639; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_640; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_641; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_642; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_643; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_644; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_645; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_646; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_647; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_648; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_649; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_650; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_651; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_652; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_653; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_654; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_655; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_656; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_657; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_658; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_659; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_660; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_661; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_662; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_663; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_664; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_665; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_666; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_667; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_668; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_669; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_670; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_671; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_672; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_673; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_674; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_675; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_676; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_677; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_678; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_679; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_680; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_681; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_682; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_683; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_684; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_685; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_686; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_687; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_688; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_689; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_690; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_691; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_692; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_693; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_694; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_695; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_696; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_697; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_698; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_699; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_700; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_701; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_702; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_703; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_704; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_705; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_706; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_707; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_708; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_709; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_710; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_711; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_712; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_713; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_714; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_715; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_716; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_717; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_718; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_719; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_720; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_721; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_722; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_723; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_724; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_725; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_726; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_727; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_728; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_729; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_730; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_731; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_732; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_733; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_734; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_735; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_736; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_737; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_738; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_739; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_740; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_741; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_742; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_743; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_744; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_745; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_746; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_747; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_748; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_749; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_750; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_751; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_752; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_753; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_754; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_755; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_756; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_757; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_758; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_759; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_760; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_761; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_762; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_763; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_764; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_765; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_766; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_767; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_768; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_769; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_770; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_771; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_772; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_773; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_774; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_775; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_776; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_777; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_778; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_779; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_780; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_781; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_782; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_783; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_784; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_785; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_786; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_787; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_788; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_789; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_790; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_791; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_792; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_793; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_794; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_795; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_796; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_797; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_798; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_799; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_800; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_801; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_802; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_803; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_804; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_805; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_806; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_807; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_808; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_809; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_810; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_811; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_812; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_813; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_814; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_815; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_816; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_817; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_818; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_819; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_820; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_821; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_822; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_823; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_824; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_825; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_826; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_827; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_828; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_829; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_830; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_831; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_832; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_833; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_834; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_835; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_836; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_837; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_838; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_839; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_840; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_841; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_842; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_843; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_844; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_845; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_846; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_847; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_848; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_849; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_850; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_851; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_852; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_853; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_854; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_855; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_856; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_857; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_858; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_859; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_860; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_861; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_862; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_863; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_864; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_865; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_866; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_867; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_868; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_869; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_870; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_871; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_872; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_873; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_874; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_875; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_876; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_877; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_878; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_879; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_880; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_881; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_882; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_883; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_884; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_885; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_886; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_887; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_888; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_889; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_890; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_891; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_892; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_893; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_894; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_895; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_896; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_897; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_898; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_899; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_900; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_901; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_902; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_903; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_904; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_905; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_906; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_907; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_908; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_909; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_910; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_911; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_912; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_913; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_914; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_915; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_916; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_917; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_918; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_919; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_920; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_921; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_922; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_923; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_924; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_925; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_926; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_927; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_928; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_929; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_930; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_931; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_932; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_933; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_934; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_935; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_936; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_937; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_938; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_939; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_940; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_941; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_942; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_943; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_944; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_945; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_946; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_947; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_948; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_949; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_950; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_951; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_952; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_953; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_954; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_955; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_956; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_957; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_958; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_959; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_960; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_961; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_962; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_963; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_964; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_965; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_966; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_967; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_968; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_969; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_970; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_971; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_972; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_973; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_974; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_975; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_976; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_977; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_978; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_979; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_980; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_981; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_982; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_983; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_984; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_985; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_986; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_987; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_988; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_989; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_990; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_991; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_992; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_993; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_994; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_995; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_996; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_997; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_998; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_999; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1000; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1001; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1002; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1003; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1004; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1005; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1006; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1007; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1008; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1009; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1010; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1011; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1012; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1013; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1014; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1015; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1016; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1017; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1018; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1019; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1020; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1021; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1022; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1023; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1024; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1025; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1026; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1027; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1028; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1029; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1030; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1031; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1032; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1033; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1034; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1035; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1036; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1037; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1038; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1039; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1040; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1041; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1042; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1043; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1044; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1045; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1046; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1047; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1048; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1049; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1050; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1051; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1052; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1053; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1054; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1055; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1056; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1057; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1058; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1059; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1060; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1061; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1062; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1063; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1064; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1065; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1066; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1067; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1068; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1069; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1070; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1071; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1072; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1073; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1074; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1075; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1076; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1077; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1078; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1079; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1080; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1081; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1082; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1083; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1084; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1085; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1086; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1087; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1088; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1089; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1090; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1091; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1092; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1093; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1094; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1095; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1096; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1097; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1098; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1099; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1100; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1101; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1102; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1103; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1104; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1105; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1106; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1107; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1108; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1109; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1110; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1111; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1112; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1113; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1114; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1115; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1116; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1117; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1118; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1119; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1120; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1121; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1122; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1123; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1124; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1125; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1126; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1127; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1128; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1129; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1130; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1131; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1132; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1133; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1134; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1135; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1136; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1137; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1138; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1139; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1140; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1141; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1142; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1143; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1144; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1145; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1146; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1147; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1148; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1149; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1150; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1151; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1152; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1153; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1154; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1155; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1156; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1157; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1158; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1159; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1160; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1161; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1162; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1163; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1164; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1165; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1166; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1167; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1168; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1169; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1170; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1171; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1172; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1173; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1174; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1175; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1176; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1177; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1178; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1179; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1180; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1181; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1182; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1183; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1184; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1185; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1186; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1187; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1188; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1189; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1190; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1191; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1192; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1193; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1194; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1195; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1196; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1197; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1198; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1199; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1200; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1201; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1202; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1203; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1204; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1205; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1206; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1207; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1208; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1209; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1210; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1211; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1212; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1213; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1214; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1215; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1216; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1217; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1218; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1219; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1220; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1221; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1222; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1223; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1224; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1225; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1226; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1227; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1228; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1229; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1230; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1231; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1232; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1233; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1234; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1235; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1236; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1237; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1238; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1239; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1240; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1241; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1242; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1243; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1244; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1245; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1246; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1247; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1248; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1249; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1250; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1251; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1252; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1253; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1254; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1255; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1256; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1257; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1258; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1259; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1260; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1261; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1262; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1263; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1264; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1265; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1266; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1267; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1268; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1269; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1270; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1271; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1272; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1273; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1274; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1275; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1276; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1277; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1278; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1279; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1280; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1281; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1282; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1283; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1284; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1285; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1286; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1287; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1288; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1289; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1290; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1291; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1292; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1293; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1294; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1295; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1296; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1297; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1298; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1299; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1300; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1301; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1302; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1303; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1304; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1305; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1306; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1307; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1308; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1309; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1310; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1311; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1312; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1313; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1314; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1315; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1316; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1317; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1318; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1319; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1320; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1321; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1322; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1323; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1324; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1325; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1326; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1327; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1328; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1329; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1330; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1331; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1332; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1333; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1334; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1335; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1336; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1337; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1338; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1339; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1340; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1341; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1342; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1343; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1344; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1345; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1346; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1347; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1348; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1349; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1350; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1351; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1352; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1353; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1354; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1355; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1356; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1357; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1358; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1359; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1360; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1361; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1362; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1363; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1364; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1365; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1366; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1367; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1368; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1369; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1370; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1371; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1372; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1373; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1374; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1375; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1376; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1377; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1378; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1379; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1380; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1381; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1382; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1383; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1384; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1385; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1386; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1387; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1388; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1389; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1390; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1391; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1392; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1393; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1394; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1395; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1396; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1397; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1398; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1399; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1400; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1401; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1402; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1403; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1404; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1405; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1406; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1407; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1408; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1409; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1410; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1411; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1412; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1413; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1414; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1415; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1416; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1417; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1418; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1419; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1420; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1421; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1422; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1423; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1424; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1425; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1426; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1427; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1428; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1429; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1430; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1431; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1432; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1433; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1434; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1435; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1436; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1437; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1438; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1439; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1440; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1441; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1442; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1443; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1444; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1445; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1446; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1447; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1448; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1449; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1450; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1451; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1452; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1453; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1454; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1455; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1456; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1457; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1458; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1459; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1460; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1461; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1462; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1463; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1464; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1465; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1466; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1467; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1468; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1469; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1470; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1471; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1472; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1473; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1474; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1475; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1476; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1477; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1478; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1479; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1480; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1481; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1482; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1483; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1484; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1485; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1486; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1487; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1488; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1489; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1490; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1491; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1492; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1493; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1494; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1495; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1496; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1497; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1498; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1499; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1500; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1501; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1502; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1503; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1504; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1505; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1506; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1507; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1508; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1509; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1510; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1511; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1512; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1513; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1514; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1515; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1516; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1517; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1518; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1519; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1520; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1521; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1522; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1523; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1524; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1525; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1526; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1527; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1528; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1529; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1530; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1531; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1532; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1533; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1534; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1535; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1536; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1537; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1538; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1539; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1540; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1541; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1542; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1543; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1544; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1545; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1546; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1547; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1548; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1549; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1550; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1551; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1552; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1553; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1554; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1555; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1556; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1557; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1558; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1559; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1560; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1561; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1562; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1563; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1564; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1565; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1566; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1567; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1568; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1569; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1570; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1571; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1572; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1573; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1574; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1575; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1576; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1577; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1578; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1579; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1580; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1581; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1582; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1583; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1584; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1585; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1586; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1587; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1588; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1589; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1590; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1591; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1592; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1593; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1594; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1595; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1596; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1597; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1598; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1599; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1600; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1601; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1602; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1603; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1604; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1605; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1606; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1607; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1608; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1609; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1610; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1611; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1612; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1613; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1614; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1615; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1616; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1617; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1618; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1619; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1620; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1621; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1622; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1623; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1624; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1625; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1626; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1627; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1628; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1629; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1630; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1631; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1632; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1633; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1634; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1635; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1636; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1637; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1638; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1639; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1640; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1641; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1642; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1643; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1644; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1645; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1646; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1647; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1648; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1649; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1650; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1651; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1652; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1653; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1654; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1655; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1656; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1657; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1658; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1659; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1660; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1661; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1662; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1663; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1664; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1665; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1666; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1667; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1668; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1669; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1670; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1671; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1672; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1673; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1674; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1675; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1676; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1677; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1678; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1679; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1680; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1681; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1682; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1683; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1684; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1685; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1686; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1687; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1688; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1689; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1690; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1691; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1692; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1693; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1694; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1695; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1696; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1697; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1698; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1699; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1700; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1701; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1702; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1703; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1704; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1705; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1706; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1707; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1708; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1709; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1710; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1711; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1712; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1713; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1714; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1715; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1716; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1717; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1718; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1719; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1720; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1721; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1722; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1723; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1724; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1725; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1726; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1727; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1728; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1729; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1730; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1731; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1732; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1733; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1734; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1735; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1736; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1737; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1738; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1739; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1740; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1741; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1742; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1743; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1744; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1745; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1746; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1747; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1748; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1749; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1750; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1751; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1752; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1753; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1754; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1755; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1756; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1757; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1758; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1759; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1760; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1761; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1762; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1763; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1764; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1765; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1766; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1767; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1768; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1769; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1770; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1771; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1772; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1773; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1774; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1775; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1776; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1777; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1778; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1779; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1780; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1781; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1782; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1783; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1784; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1785; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1786; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1787; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1788; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1789; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1790; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1791; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1792; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1793; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1794; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1795; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1796; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1797; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1798; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1799; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1800; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1801; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1802; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1803; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1804; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1805; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1806; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1807; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1808; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1809; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1810; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1811; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1812; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1813; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1814; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1815; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1816; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1817; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1818; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1819; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1820; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1821; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1822; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1823; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1824; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1825; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1826; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1827; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1828; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1829; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1830; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1831; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1832; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1833; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1834; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1835; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1836; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1837; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1838; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1839; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1840; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1841; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1842; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1843; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1844; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1845; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1846; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1847; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1848; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1849; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1850; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1851; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1852; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1853; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1854; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1855; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1856; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1857; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1858; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1859; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1860; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1861; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1862; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1863; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1864; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1865; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1866; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1867; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1868; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1869; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1870; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1871; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1872; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1873; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1874; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1875; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1876; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1877; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1878; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1879; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1880; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1881; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1882; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1883; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1884; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1885; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1886; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1887; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1888; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1889; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1890; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1891; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1892; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1893; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1894; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1895; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1896; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1897; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1898; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1899; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1900; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1901; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1902; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1903; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1904; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1905; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1906; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1907; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1908; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1909; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1910; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1911; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1912; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1913; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1914; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1915; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1916; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1917; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1918; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1919; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1920; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1921; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1922; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1923; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1924; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1925; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1926; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1927; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1928; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1929; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1930; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1931; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1932; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1933; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1934; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1935; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1936; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1937; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1938; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1939; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1940; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1941; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1942; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1943; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1944; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1945; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1946; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1947; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1948; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1949; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1950; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1951; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1952; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1953; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1954; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1955; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1956; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1957; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1958; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1959; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1960; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1961; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1962; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1963; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1964; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1965; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1966; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1967; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1968; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1969; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1970; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1971; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1972; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1973; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1974; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1975; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1976; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1977; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1978; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1979; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1980; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1981; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1982; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1983; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1984; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1985; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1986; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1987; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1988; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1989; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1990; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1991; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1992; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1993; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1994; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1995; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1996; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1997; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1998; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_1999; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_2000; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_2001; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_2002; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_2003; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_2004; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_2005; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_2006; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_2007; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_2008; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_2009; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_2010; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_2011; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_2012; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_2013; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_2014; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_2015; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_2016; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_2017; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_2018; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_2019; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_2020; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_2021; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_2022; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_2023; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_2024; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_2025; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_2026; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_2027; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_2028; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_2029; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_2030; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_2031; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_2032; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_2033; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_2034; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_2035; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_2036; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_2037; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_2038; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_2039; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_2040; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_2041; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_2042; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_2043; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_2044; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_2045; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_2046; // @[Multiplier.scala 64:55]
  wire [9:0] _GEN_2047; // @[Multiplier.scala 64:55]
  wire [9:0] _T_10; // @[Multiplier.scala 64:55]
  wire [8:0] _T_11; // @[Multiplier.scala 64:100]
  wire [520:0] _GEN_2048; // @[Multiplier.scala 64:91]
  wire [520:0] _T_12; // @[Multiplier.scala 64:91]
  wire  _T_13; // @[Multiplier.scala 66:34]
  wire [5:0] _T_16; // @[Multiplier.scala 66:57]
  wire [8:0] _GEN_2049; // @[Multiplier.scala 66:55]
  wire  _T_17; // @[Multiplier.scala 66:55]
  wire  _T_19; // @[Multiplier.scala 67:32]
  wire  _T_20; // @[Multiplier.scala 67:52]
  wire  _T_22; // @[Multiplier.scala 68:42]
  wire  _T_23; // @[Multiplier.scala 68:76]
  wire [520:0] _T_25; // @[Multiplier.scala 68:105]
  wire [520:0] _T_28; // @[Multiplier.scala 68:97]
  wire [520:0] _T_30; // @[Multiplier.scala 68:64]
  wire [520:0] _T_31; // @[Multiplier.scala 68:29]
  assign exponentSum = $signed(io_A_exponent) + $signed(io_B_exponent); // @[Multiplier.scala 60:49]
  assign fractionSum = io_A_fraction[11:0] + io_B_fraction[11:0]; // @[Multiplier.scala 61:71]
  assign _T_4 = 7'sh38 + $signed(exponentSum); // @[Multiplier.scala 63:42]
  assign shift = $signed(_T_4) - 8'sh8; // @[Multiplier.scala 63:57]
  assign _T_5 = $signed(shift) < 9'sh0; // @[Multiplier.scala 64:32]
  assign _T_9 = 9'sh0 - $signed(shift); // @[Multiplier.scala 64:67]
  assign _GEN_3 = 11'h3 == fractionSum[12:2] ? 10'h101 : 10'h100; // @[Multiplier.scala 64:55]
  assign _GEN_4 = 11'h4 == fractionSum[12:2] ? 10'h101 : _GEN_3; // @[Multiplier.scala 64:55]
  assign _GEN_5 = 11'h5 == fractionSum[12:2] ? 10'h101 : _GEN_4; // @[Multiplier.scala 64:55]
  assign _GEN_6 = 11'h6 == fractionSum[12:2] ? 10'h101 : _GEN_5; // @[Multiplier.scala 64:55]
  assign _GEN_7 = 11'h7 == fractionSum[12:2] ? 10'h101 : _GEN_6; // @[Multiplier.scala 64:55]
  assign _GEN_8 = 11'h8 == fractionSum[12:2] ? 10'h101 : _GEN_7; // @[Multiplier.scala 64:55]
  assign _GEN_9 = 11'h9 == fractionSum[12:2] ? 10'h102 : _GEN_8; // @[Multiplier.scala 64:55]
  assign _GEN_10 = 11'ha == fractionSum[12:2] ? 10'h102 : _GEN_9; // @[Multiplier.scala 64:55]
  assign _GEN_11 = 11'hb == fractionSum[12:2] ? 10'h102 : _GEN_10; // @[Multiplier.scala 64:55]
  assign _GEN_12 = 11'hc == fractionSum[12:2] ? 10'h102 : _GEN_11; // @[Multiplier.scala 64:55]
  assign _GEN_13 = 11'hd == fractionSum[12:2] ? 10'h102 : _GEN_12; // @[Multiplier.scala 64:55]
  assign _GEN_14 = 11'he == fractionSum[12:2] ? 10'h102 : _GEN_13; // @[Multiplier.scala 64:55]
  assign _GEN_15 = 11'hf == fractionSum[12:2] ? 10'h103 : _GEN_14; // @[Multiplier.scala 64:55]
  assign _GEN_16 = 11'h10 == fractionSum[12:2] ? 10'h103 : _GEN_15; // @[Multiplier.scala 64:55]
  assign _GEN_17 = 11'h11 == fractionSum[12:2] ? 10'h103 : _GEN_16; // @[Multiplier.scala 64:55]
  assign _GEN_18 = 11'h12 == fractionSum[12:2] ? 10'h103 : _GEN_17; // @[Multiplier.scala 64:55]
  assign _GEN_19 = 11'h13 == fractionSum[12:2] ? 10'h103 : _GEN_18; // @[Multiplier.scala 64:55]
  assign _GEN_20 = 11'h14 == fractionSum[12:2] ? 10'h103 : _GEN_19; // @[Multiplier.scala 64:55]
  assign _GEN_21 = 11'h15 == fractionSum[12:2] ? 10'h104 : _GEN_20; // @[Multiplier.scala 64:55]
  assign _GEN_22 = 11'h16 == fractionSum[12:2] ? 10'h104 : _GEN_21; // @[Multiplier.scala 64:55]
  assign _GEN_23 = 11'h17 == fractionSum[12:2] ? 10'h104 : _GEN_22; // @[Multiplier.scala 64:55]
  assign _GEN_24 = 11'h18 == fractionSum[12:2] ? 10'h104 : _GEN_23; // @[Multiplier.scala 64:55]
  assign _GEN_25 = 11'h19 == fractionSum[12:2] ? 10'h104 : _GEN_24; // @[Multiplier.scala 64:55]
  assign _GEN_26 = 11'h1a == fractionSum[12:2] ? 10'h105 : _GEN_25; // @[Multiplier.scala 64:55]
  assign _GEN_27 = 11'h1b == fractionSum[12:2] ? 10'h105 : _GEN_26; // @[Multiplier.scala 64:55]
  assign _GEN_28 = 11'h1c == fractionSum[12:2] ? 10'h105 : _GEN_27; // @[Multiplier.scala 64:55]
  assign _GEN_29 = 11'h1d == fractionSum[12:2] ? 10'h105 : _GEN_28; // @[Multiplier.scala 64:55]
  assign _GEN_30 = 11'h1e == fractionSum[12:2] ? 10'h105 : _GEN_29; // @[Multiplier.scala 64:55]
  assign _GEN_31 = 11'h1f == fractionSum[12:2] ? 10'h105 : _GEN_30; // @[Multiplier.scala 64:55]
  assign _GEN_32 = 11'h20 == fractionSum[12:2] ? 10'h106 : _GEN_31; // @[Multiplier.scala 64:55]
  assign _GEN_33 = 11'h21 == fractionSum[12:2] ? 10'h106 : _GEN_32; // @[Multiplier.scala 64:55]
  assign _GEN_34 = 11'h22 == fractionSum[12:2] ? 10'h106 : _GEN_33; // @[Multiplier.scala 64:55]
  assign _GEN_35 = 11'h23 == fractionSum[12:2] ? 10'h106 : _GEN_34; // @[Multiplier.scala 64:55]
  assign _GEN_36 = 11'h24 == fractionSum[12:2] ? 10'h106 : _GEN_35; // @[Multiplier.scala 64:55]
  assign _GEN_37 = 11'h25 == fractionSum[12:2] ? 10'h106 : _GEN_36; // @[Multiplier.scala 64:55]
  assign _GEN_38 = 11'h26 == fractionSum[12:2] ? 10'h107 : _GEN_37; // @[Multiplier.scala 64:55]
  assign _GEN_39 = 11'h27 == fractionSum[12:2] ? 10'h107 : _GEN_38; // @[Multiplier.scala 64:55]
  assign _GEN_40 = 11'h28 == fractionSum[12:2] ? 10'h107 : _GEN_39; // @[Multiplier.scala 64:55]
  assign _GEN_41 = 11'h29 == fractionSum[12:2] ? 10'h107 : _GEN_40; // @[Multiplier.scala 64:55]
  assign _GEN_42 = 11'h2a == fractionSum[12:2] ? 10'h107 : _GEN_41; // @[Multiplier.scala 64:55]
  assign _GEN_43 = 11'h2b == fractionSum[12:2] ? 10'h108 : _GEN_42; // @[Multiplier.scala 64:55]
  assign _GEN_44 = 11'h2c == fractionSum[12:2] ? 10'h108 : _GEN_43; // @[Multiplier.scala 64:55]
  assign _GEN_45 = 11'h2d == fractionSum[12:2] ? 10'h108 : _GEN_44; // @[Multiplier.scala 64:55]
  assign _GEN_46 = 11'h2e == fractionSum[12:2] ? 10'h108 : _GEN_45; // @[Multiplier.scala 64:55]
  assign _GEN_47 = 11'h2f == fractionSum[12:2] ? 10'h108 : _GEN_46; // @[Multiplier.scala 64:55]
  assign _GEN_48 = 11'h30 == fractionSum[12:2] ? 10'h108 : _GEN_47; // @[Multiplier.scala 64:55]
  assign _GEN_49 = 11'h31 == fractionSum[12:2] ? 10'h109 : _GEN_48; // @[Multiplier.scala 64:55]
  assign _GEN_50 = 11'h32 == fractionSum[12:2] ? 10'h109 : _GEN_49; // @[Multiplier.scala 64:55]
  assign _GEN_51 = 11'h33 == fractionSum[12:2] ? 10'h109 : _GEN_50; // @[Multiplier.scala 64:55]
  assign _GEN_52 = 11'h34 == fractionSum[12:2] ? 10'h109 : _GEN_51; // @[Multiplier.scala 64:55]
  assign _GEN_53 = 11'h35 == fractionSum[12:2] ? 10'h109 : _GEN_52; // @[Multiplier.scala 64:55]
  assign _GEN_54 = 11'h36 == fractionSum[12:2] ? 10'h10a : _GEN_53; // @[Multiplier.scala 64:55]
  assign _GEN_55 = 11'h37 == fractionSum[12:2] ? 10'h10a : _GEN_54; // @[Multiplier.scala 64:55]
  assign _GEN_56 = 11'h38 == fractionSum[12:2] ? 10'h10a : _GEN_55; // @[Multiplier.scala 64:55]
  assign _GEN_57 = 11'h39 == fractionSum[12:2] ? 10'h10a : _GEN_56; // @[Multiplier.scala 64:55]
  assign _GEN_58 = 11'h3a == fractionSum[12:2] ? 10'h10a : _GEN_57; // @[Multiplier.scala 64:55]
  assign _GEN_59 = 11'h3b == fractionSum[12:2] ? 10'h10a : _GEN_58; // @[Multiplier.scala 64:55]
  assign _GEN_60 = 11'h3c == fractionSum[12:2] ? 10'h10b : _GEN_59; // @[Multiplier.scala 64:55]
  assign _GEN_61 = 11'h3d == fractionSum[12:2] ? 10'h10b : _GEN_60; // @[Multiplier.scala 64:55]
  assign _GEN_62 = 11'h3e == fractionSum[12:2] ? 10'h10b : _GEN_61; // @[Multiplier.scala 64:55]
  assign _GEN_63 = 11'h3f == fractionSum[12:2] ? 10'h10b : _GEN_62; // @[Multiplier.scala 64:55]
  assign _GEN_64 = 11'h40 == fractionSum[12:2] ? 10'h10b : _GEN_63; // @[Multiplier.scala 64:55]
  assign _GEN_65 = 11'h41 == fractionSum[12:2] ? 10'h10c : _GEN_64; // @[Multiplier.scala 64:55]
  assign _GEN_66 = 11'h42 == fractionSum[12:2] ? 10'h10c : _GEN_65; // @[Multiplier.scala 64:55]
  assign _GEN_67 = 11'h43 == fractionSum[12:2] ? 10'h10c : _GEN_66; // @[Multiplier.scala 64:55]
  assign _GEN_68 = 11'h44 == fractionSum[12:2] ? 10'h10c : _GEN_67; // @[Multiplier.scala 64:55]
  assign _GEN_69 = 11'h45 == fractionSum[12:2] ? 10'h10c : _GEN_68; // @[Multiplier.scala 64:55]
  assign _GEN_70 = 11'h46 == fractionSum[12:2] ? 10'h10c : _GEN_69; // @[Multiplier.scala 64:55]
  assign _GEN_71 = 11'h47 == fractionSum[12:2] ? 10'h10d : _GEN_70; // @[Multiplier.scala 64:55]
  assign _GEN_72 = 11'h48 == fractionSum[12:2] ? 10'h10d : _GEN_71; // @[Multiplier.scala 64:55]
  assign _GEN_73 = 11'h49 == fractionSum[12:2] ? 10'h10d : _GEN_72; // @[Multiplier.scala 64:55]
  assign _GEN_74 = 11'h4a == fractionSum[12:2] ? 10'h10d : _GEN_73; // @[Multiplier.scala 64:55]
  assign _GEN_75 = 11'h4b == fractionSum[12:2] ? 10'h10d : _GEN_74; // @[Multiplier.scala 64:55]
  assign _GEN_76 = 11'h4c == fractionSum[12:2] ? 10'h10e : _GEN_75; // @[Multiplier.scala 64:55]
  assign _GEN_77 = 11'h4d == fractionSum[12:2] ? 10'h10e : _GEN_76; // @[Multiplier.scala 64:55]
  assign _GEN_78 = 11'h4e == fractionSum[12:2] ? 10'h10e : _GEN_77; // @[Multiplier.scala 64:55]
  assign _GEN_79 = 11'h4f == fractionSum[12:2] ? 10'h10e : _GEN_78; // @[Multiplier.scala 64:55]
  assign _GEN_80 = 11'h50 == fractionSum[12:2] ? 10'h10e : _GEN_79; // @[Multiplier.scala 64:55]
  assign _GEN_81 = 11'h51 == fractionSum[12:2] ? 10'h10e : _GEN_80; // @[Multiplier.scala 64:55]
  assign _GEN_82 = 11'h52 == fractionSum[12:2] ? 10'h10f : _GEN_81; // @[Multiplier.scala 64:55]
  assign _GEN_83 = 11'h53 == fractionSum[12:2] ? 10'h10f : _GEN_82; // @[Multiplier.scala 64:55]
  assign _GEN_84 = 11'h54 == fractionSum[12:2] ? 10'h10f : _GEN_83; // @[Multiplier.scala 64:55]
  assign _GEN_85 = 11'h55 == fractionSum[12:2] ? 10'h10f : _GEN_84; // @[Multiplier.scala 64:55]
  assign _GEN_86 = 11'h56 == fractionSum[12:2] ? 10'h10f : _GEN_85; // @[Multiplier.scala 64:55]
  assign _GEN_87 = 11'h57 == fractionSum[12:2] ? 10'h110 : _GEN_86; // @[Multiplier.scala 64:55]
  assign _GEN_88 = 11'h58 == fractionSum[12:2] ? 10'h110 : _GEN_87; // @[Multiplier.scala 64:55]
  assign _GEN_89 = 11'h59 == fractionSum[12:2] ? 10'h110 : _GEN_88; // @[Multiplier.scala 64:55]
  assign _GEN_90 = 11'h5a == fractionSum[12:2] ? 10'h110 : _GEN_89; // @[Multiplier.scala 64:55]
  assign _GEN_91 = 11'h5b == fractionSum[12:2] ? 10'h110 : _GEN_90; // @[Multiplier.scala 64:55]
  assign _GEN_92 = 11'h5c == fractionSum[12:2] ? 10'h110 : _GEN_91; // @[Multiplier.scala 64:55]
  assign _GEN_93 = 11'h5d == fractionSum[12:2] ? 10'h111 : _GEN_92; // @[Multiplier.scala 64:55]
  assign _GEN_94 = 11'h5e == fractionSum[12:2] ? 10'h111 : _GEN_93; // @[Multiplier.scala 64:55]
  assign _GEN_95 = 11'h5f == fractionSum[12:2] ? 10'h111 : _GEN_94; // @[Multiplier.scala 64:55]
  assign _GEN_96 = 11'h60 == fractionSum[12:2] ? 10'h111 : _GEN_95; // @[Multiplier.scala 64:55]
  assign _GEN_97 = 11'h61 == fractionSum[12:2] ? 10'h111 : _GEN_96; // @[Multiplier.scala 64:55]
  assign _GEN_98 = 11'h62 == fractionSum[12:2] ? 10'h112 : _GEN_97; // @[Multiplier.scala 64:55]
  assign _GEN_99 = 11'h63 == fractionSum[12:2] ? 10'h112 : _GEN_98; // @[Multiplier.scala 64:55]
  assign _GEN_100 = 11'h64 == fractionSum[12:2] ? 10'h112 : _GEN_99; // @[Multiplier.scala 64:55]
  assign _GEN_101 = 11'h65 == fractionSum[12:2] ? 10'h112 : _GEN_100; // @[Multiplier.scala 64:55]
  assign _GEN_102 = 11'h66 == fractionSum[12:2] ? 10'h112 : _GEN_101; // @[Multiplier.scala 64:55]
  assign _GEN_103 = 11'h67 == fractionSum[12:2] ? 10'h112 : _GEN_102; // @[Multiplier.scala 64:55]
  assign _GEN_104 = 11'h68 == fractionSum[12:2] ? 10'h113 : _GEN_103; // @[Multiplier.scala 64:55]
  assign _GEN_105 = 11'h69 == fractionSum[12:2] ? 10'h113 : _GEN_104; // @[Multiplier.scala 64:55]
  assign _GEN_106 = 11'h6a == fractionSum[12:2] ? 10'h113 : _GEN_105; // @[Multiplier.scala 64:55]
  assign _GEN_107 = 11'h6b == fractionSum[12:2] ? 10'h113 : _GEN_106; // @[Multiplier.scala 64:55]
  assign _GEN_108 = 11'h6c == fractionSum[12:2] ? 10'h113 : _GEN_107; // @[Multiplier.scala 64:55]
  assign _GEN_109 = 11'h6d == fractionSum[12:2] ? 10'h114 : _GEN_108; // @[Multiplier.scala 64:55]
  assign _GEN_110 = 11'h6e == fractionSum[12:2] ? 10'h114 : _GEN_109; // @[Multiplier.scala 64:55]
  assign _GEN_111 = 11'h6f == fractionSum[12:2] ? 10'h114 : _GEN_110; // @[Multiplier.scala 64:55]
  assign _GEN_112 = 11'h70 == fractionSum[12:2] ? 10'h114 : _GEN_111; // @[Multiplier.scala 64:55]
  assign _GEN_113 = 11'h71 == fractionSum[12:2] ? 10'h114 : _GEN_112; // @[Multiplier.scala 64:55]
  assign _GEN_114 = 11'h72 == fractionSum[12:2] ? 10'h115 : _GEN_113; // @[Multiplier.scala 64:55]
  assign _GEN_115 = 11'h73 == fractionSum[12:2] ? 10'h115 : _GEN_114; // @[Multiplier.scala 64:55]
  assign _GEN_116 = 11'h74 == fractionSum[12:2] ? 10'h115 : _GEN_115; // @[Multiplier.scala 64:55]
  assign _GEN_117 = 11'h75 == fractionSum[12:2] ? 10'h115 : _GEN_116; // @[Multiplier.scala 64:55]
  assign _GEN_118 = 11'h76 == fractionSum[12:2] ? 10'h115 : _GEN_117; // @[Multiplier.scala 64:55]
  assign _GEN_119 = 11'h77 == fractionSum[12:2] ? 10'h115 : _GEN_118; // @[Multiplier.scala 64:55]
  assign _GEN_120 = 11'h78 == fractionSum[12:2] ? 10'h116 : _GEN_119; // @[Multiplier.scala 64:55]
  assign _GEN_121 = 11'h79 == fractionSum[12:2] ? 10'h116 : _GEN_120; // @[Multiplier.scala 64:55]
  assign _GEN_122 = 11'h7a == fractionSum[12:2] ? 10'h116 : _GEN_121; // @[Multiplier.scala 64:55]
  assign _GEN_123 = 11'h7b == fractionSum[12:2] ? 10'h116 : _GEN_122; // @[Multiplier.scala 64:55]
  assign _GEN_124 = 11'h7c == fractionSum[12:2] ? 10'h116 : _GEN_123; // @[Multiplier.scala 64:55]
  assign _GEN_125 = 11'h7d == fractionSum[12:2] ? 10'h117 : _GEN_124; // @[Multiplier.scala 64:55]
  assign _GEN_126 = 11'h7e == fractionSum[12:2] ? 10'h117 : _GEN_125; // @[Multiplier.scala 64:55]
  assign _GEN_127 = 11'h7f == fractionSum[12:2] ? 10'h117 : _GEN_126; // @[Multiplier.scala 64:55]
  assign _GEN_128 = 11'h80 == fractionSum[12:2] ? 10'h117 : _GEN_127; // @[Multiplier.scala 64:55]
  assign _GEN_129 = 11'h81 == fractionSum[12:2] ? 10'h117 : _GEN_128; // @[Multiplier.scala 64:55]
  assign _GEN_130 = 11'h82 == fractionSum[12:2] ? 10'h118 : _GEN_129; // @[Multiplier.scala 64:55]
  assign _GEN_131 = 11'h83 == fractionSum[12:2] ? 10'h118 : _GEN_130; // @[Multiplier.scala 64:55]
  assign _GEN_132 = 11'h84 == fractionSum[12:2] ? 10'h118 : _GEN_131; // @[Multiplier.scala 64:55]
  assign _GEN_133 = 11'h85 == fractionSum[12:2] ? 10'h118 : _GEN_132; // @[Multiplier.scala 64:55]
  assign _GEN_134 = 11'h86 == fractionSum[12:2] ? 10'h118 : _GEN_133; // @[Multiplier.scala 64:55]
  assign _GEN_135 = 11'h87 == fractionSum[12:2] ? 10'h118 : _GEN_134; // @[Multiplier.scala 64:55]
  assign _GEN_136 = 11'h88 == fractionSum[12:2] ? 10'h119 : _GEN_135; // @[Multiplier.scala 64:55]
  assign _GEN_137 = 11'h89 == fractionSum[12:2] ? 10'h119 : _GEN_136; // @[Multiplier.scala 64:55]
  assign _GEN_138 = 11'h8a == fractionSum[12:2] ? 10'h119 : _GEN_137; // @[Multiplier.scala 64:55]
  assign _GEN_139 = 11'h8b == fractionSum[12:2] ? 10'h119 : _GEN_138; // @[Multiplier.scala 64:55]
  assign _GEN_140 = 11'h8c == fractionSum[12:2] ? 10'h119 : _GEN_139; // @[Multiplier.scala 64:55]
  assign _GEN_141 = 11'h8d == fractionSum[12:2] ? 10'h11a : _GEN_140; // @[Multiplier.scala 64:55]
  assign _GEN_142 = 11'h8e == fractionSum[12:2] ? 10'h11a : _GEN_141; // @[Multiplier.scala 64:55]
  assign _GEN_143 = 11'h8f == fractionSum[12:2] ? 10'h11a : _GEN_142; // @[Multiplier.scala 64:55]
  assign _GEN_144 = 11'h90 == fractionSum[12:2] ? 10'h11a : _GEN_143; // @[Multiplier.scala 64:55]
  assign _GEN_145 = 11'h91 == fractionSum[12:2] ? 10'h11a : _GEN_144; // @[Multiplier.scala 64:55]
  assign _GEN_146 = 11'h92 == fractionSum[12:2] ? 10'h11b : _GEN_145; // @[Multiplier.scala 64:55]
  assign _GEN_147 = 11'h93 == fractionSum[12:2] ? 10'h11b : _GEN_146; // @[Multiplier.scala 64:55]
  assign _GEN_148 = 11'h94 == fractionSum[12:2] ? 10'h11b : _GEN_147; // @[Multiplier.scala 64:55]
  assign _GEN_149 = 11'h95 == fractionSum[12:2] ? 10'h11b : _GEN_148; // @[Multiplier.scala 64:55]
  assign _GEN_150 = 11'h96 == fractionSum[12:2] ? 10'h11b : _GEN_149; // @[Multiplier.scala 64:55]
  assign _GEN_151 = 11'h97 == fractionSum[12:2] ? 10'h11c : _GEN_150; // @[Multiplier.scala 64:55]
  assign _GEN_152 = 11'h98 == fractionSum[12:2] ? 10'h11c : _GEN_151; // @[Multiplier.scala 64:55]
  assign _GEN_153 = 11'h99 == fractionSum[12:2] ? 10'h11c : _GEN_152; // @[Multiplier.scala 64:55]
  assign _GEN_154 = 11'h9a == fractionSum[12:2] ? 10'h11c : _GEN_153; // @[Multiplier.scala 64:55]
  assign _GEN_155 = 11'h9b == fractionSum[12:2] ? 10'h11c : _GEN_154; // @[Multiplier.scala 64:55]
  assign _GEN_156 = 11'h9c == fractionSum[12:2] ? 10'h11d : _GEN_155; // @[Multiplier.scala 64:55]
  assign _GEN_157 = 11'h9d == fractionSum[12:2] ? 10'h11d : _GEN_156; // @[Multiplier.scala 64:55]
  assign _GEN_158 = 11'h9e == fractionSum[12:2] ? 10'h11d : _GEN_157; // @[Multiplier.scala 64:55]
  assign _GEN_159 = 11'h9f == fractionSum[12:2] ? 10'h11d : _GEN_158; // @[Multiplier.scala 64:55]
  assign _GEN_160 = 11'ha0 == fractionSum[12:2] ? 10'h11d : _GEN_159; // @[Multiplier.scala 64:55]
  assign _GEN_161 = 11'ha1 == fractionSum[12:2] ? 10'h11d : _GEN_160; // @[Multiplier.scala 64:55]
  assign _GEN_162 = 11'ha2 == fractionSum[12:2] ? 10'h11e : _GEN_161; // @[Multiplier.scala 64:55]
  assign _GEN_163 = 11'ha3 == fractionSum[12:2] ? 10'h11e : _GEN_162; // @[Multiplier.scala 64:55]
  assign _GEN_164 = 11'ha4 == fractionSum[12:2] ? 10'h11e : _GEN_163; // @[Multiplier.scala 64:55]
  assign _GEN_165 = 11'ha5 == fractionSum[12:2] ? 10'h11e : _GEN_164; // @[Multiplier.scala 64:55]
  assign _GEN_166 = 11'ha6 == fractionSum[12:2] ? 10'h11e : _GEN_165; // @[Multiplier.scala 64:55]
  assign _GEN_167 = 11'ha7 == fractionSum[12:2] ? 10'h11f : _GEN_166; // @[Multiplier.scala 64:55]
  assign _GEN_168 = 11'ha8 == fractionSum[12:2] ? 10'h11f : _GEN_167; // @[Multiplier.scala 64:55]
  assign _GEN_169 = 11'ha9 == fractionSum[12:2] ? 10'h11f : _GEN_168; // @[Multiplier.scala 64:55]
  assign _GEN_170 = 11'haa == fractionSum[12:2] ? 10'h11f : _GEN_169; // @[Multiplier.scala 64:55]
  assign _GEN_171 = 11'hab == fractionSum[12:2] ? 10'h11f : _GEN_170; // @[Multiplier.scala 64:55]
  assign _GEN_172 = 11'hac == fractionSum[12:2] ? 10'h120 : _GEN_171; // @[Multiplier.scala 64:55]
  assign _GEN_173 = 11'had == fractionSum[12:2] ? 10'h120 : _GEN_172; // @[Multiplier.scala 64:55]
  assign _GEN_174 = 11'hae == fractionSum[12:2] ? 10'h120 : _GEN_173; // @[Multiplier.scala 64:55]
  assign _GEN_175 = 11'haf == fractionSum[12:2] ? 10'h120 : _GEN_174; // @[Multiplier.scala 64:55]
  assign _GEN_176 = 11'hb0 == fractionSum[12:2] ? 10'h120 : _GEN_175; // @[Multiplier.scala 64:55]
  assign _GEN_177 = 11'hb1 == fractionSum[12:2] ? 10'h121 : _GEN_176; // @[Multiplier.scala 64:55]
  assign _GEN_178 = 11'hb2 == fractionSum[12:2] ? 10'h121 : _GEN_177; // @[Multiplier.scala 64:55]
  assign _GEN_179 = 11'hb3 == fractionSum[12:2] ? 10'h121 : _GEN_178; // @[Multiplier.scala 64:55]
  assign _GEN_180 = 11'hb4 == fractionSum[12:2] ? 10'h121 : _GEN_179; // @[Multiplier.scala 64:55]
  assign _GEN_181 = 11'hb5 == fractionSum[12:2] ? 10'h121 : _GEN_180; // @[Multiplier.scala 64:55]
  assign _GEN_182 = 11'hb6 == fractionSum[12:2] ? 10'h122 : _GEN_181; // @[Multiplier.scala 64:55]
  assign _GEN_183 = 11'hb7 == fractionSum[12:2] ? 10'h122 : _GEN_182; // @[Multiplier.scala 64:55]
  assign _GEN_184 = 11'hb8 == fractionSum[12:2] ? 10'h122 : _GEN_183; // @[Multiplier.scala 64:55]
  assign _GEN_185 = 11'hb9 == fractionSum[12:2] ? 10'h122 : _GEN_184; // @[Multiplier.scala 64:55]
  assign _GEN_186 = 11'hba == fractionSum[12:2] ? 10'h122 : _GEN_185; // @[Multiplier.scala 64:55]
  assign _GEN_187 = 11'hbb == fractionSum[12:2] ? 10'h123 : _GEN_186; // @[Multiplier.scala 64:55]
  assign _GEN_188 = 11'hbc == fractionSum[12:2] ? 10'h123 : _GEN_187; // @[Multiplier.scala 64:55]
  assign _GEN_189 = 11'hbd == fractionSum[12:2] ? 10'h123 : _GEN_188; // @[Multiplier.scala 64:55]
  assign _GEN_190 = 11'hbe == fractionSum[12:2] ? 10'h123 : _GEN_189; // @[Multiplier.scala 64:55]
  assign _GEN_191 = 11'hbf == fractionSum[12:2] ? 10'h123 : _GEN_190; // @[Multiplier.scala 64:55]
  assign _GEN_192 = 11'hc0 == fractionSum[12:2] ? 10'h124 : _GEN_191; // @[Multiplier.scala 64:55]
  assign _GEN_193 = 11'hc1 == fractionSum[12:2] ? 10'h124 : _GEN_192; // @[Multiplier.scala 64:55]
  assign _GEN_194 = 11'hc2 == fractionSum[12:2] ? 10'h124 : _GEN_193; // @[Multiplier.scala 64:55]
  assign _GEN_195 = 11'hc3 == fractionSum[12:2] ? 10'h124 : _GEN_194; // @[Multiplier.scala 64:55]
  assign _GEN_196 = 11'hc4 == fractionSum[12:2] ? 10'h124 : _GEN_195; // @[Multiplier.scala 64:55]
  assign _GEN_197 = 11'hc5 == fractionSum[12:2] ? 10'h125 : _GEN_196; // @[Multiplier.scala 64:55]
  assign _GEN_198 = 11'hc6 == fractionSum[12:2] ? 10'h125 : _GEN_197; // @[Multiplier.scala 64:55]
  assign _GEN_199 = 11'hc7 == fractionSum[12:2] ? 10'h125 : _GEN_198; // @[Multiplier.scala 64:55]
  assign _GEN_200 = 11'hc8 == fractionSum[12:2] ? 10'h125 : _GEN_199; // @[Multiplier.scala 64:55]
  assign _GEN_201 = 11'hc9 == fractionSum[12:2] ? 10'h125 : _GEN_200; // @[Multiplier.scala 64:55]
  assign _GEN_202 = 11'hca == fractionSum[12:2] ? 10'h126 : _GEN_201; // @[Multiplier.scala 64:55]
  assign _GEN_203 = 11'hcb == fractionSum[12:2] ? 10'h126 : _GEN_202; // @[Multiplier.scala 64:55]
  assign _GEN_204 = 11'hcc == fractionSum[12:2] ? 10'h126 : _GEN_203; // @[Multiplier.scala 64:55]
  assign _GEN_205 = 11'hcd == fractionSum[12:2] ? 10'h126 : _GEN_204; // @[Multiplier.scala 64:55]
  assign _GEN_206 = 11'hce == fractionSum[12:2] ? 10'h126 : _GEN_205; // @[Multiplier.scala 64:55]
  assign _GEN_207 = 11'hcf == fractionSum[12:2] ? 10'h127 : _GEN_206; // @[Multiplier.scala 64:55]
  assign _GEN_208 = 11'hd0 == fractionSum[12:2] ? 10'h127 : _GEN_207; // @[Multiplier.scala 64:55]
  assign _GEN_209 = 11'hd1 == fractionSum[12:2] ? 10'h127 : _GEN_208; // @[Multiplier.scala 64:55]
  assign _GEN_210 = 11'hd2 == fractionSum[12:2] ? 10'h127 : _GEN_209; // @[Multiplier.scala 64:55]
  assign _GEN_211 = 11'hd3 == fractionSum[12:2] ? 10'h127 : _GEN_210; // @[Multiplier.scala 64:55]
  assign _GEN_212 = 11'hd4 == fractionSum[12:2] ? 10'h128 : _GEN_211; // @[Multiplier.scala 64:55]
  assign _GEN_213 = 11'hd5 == fractionSum[12:2] ? 10'h128 : _GEN_212; // @[Multiplier.scala 64:55]
  assign _GEN_214 = 11'hd6 == fractionSum[12:2] ? 10'h128 : _GEN_213; // @[Multiplier.scala 64:55]
  assign _GEN_215 = 11'hd7 == fractionSum[12:2] ? 10'h128 : _GEN_214; // @[Multiplier.scala 64:55]
  assign _GEN_216 = 11'hd8 == fractionSum[12:2] ? 10'h128 : _GEN_215; // @[Multiplier.scala 64:55]
  assign _GEN_217 = 11'hd9 == fractionSum[12:2] ? 10'h129 : _GEN_216; // @[Multiplier.scala 64:55]
  assign _GEN_218 = 11'hda == fractionSum[12:2] ? 10'h129 : _GEN_217; // @[Multiplier.scala 64:55]
  assign _GEN_219 = 11'hdb == fractionSum[12:2] ? 10'h129 : _GEN_218; // @[Multiplier.scala 64:55]
  assign _GEN_220 = 11'hdc == fractionSum[12:2] ? 10'h129 : _GEN_219; // @[Multiplier.scala 64:55]
  assign _GEN_221 = 11'hdd == fractionSum[12:2] ? 10'h129 : _GEN_220; // @[Multiplier.scala 64:55]
  assign _GEN_222 = 11'hde == fractionSum[12:2] ? 10'h12a : _GEN_221; // @[Multiplier.scala 64:55]
  assign _GEN_223 = 11'hdf == fractionSum[12:2] ? 10'h12a : _GEN_222; // @[Multiplier.scala 64:55]
  assign _GEN_224 = 11'he0 == fractionSum[12:2] ? 10'h12a : _GEN_223; // @[Multiplier.scala 64:55]
  assign _GEN_225 = 11'he1 == fractionSum[12:2] ? 10'h12a : _GEN_224; // @[Multiplier.scala 64:55]
  assign _GEN_226 = 11'he2 == fractionSum[12:2] ? 10'h12a : _GEN_225; // @[Multiplier.scala 64:55]
  assign _GEN_227 = 11'he3 == fractionSum[12:2] ? 10'h12b : _GEN_226; // @[Multiplier.scala 64:55]
  assign _GEN_228 = 11'he4 == fractionSum[12:2] ? 10'h12b : _GEN_227; // @[Multiplier.scala 64:55]
  assign _GEN_229 = 11'he5 == fractionSum[12:2] ? 10'h12b : _GEN_228; // @[Multiplier.scala 64:55]
  assign _GEN_230 = 11'he6 == fractionSum[12:2] ? 10'h12b : _GEN_229; // @[Multiplier.scala 64:55]
  assign _GEN_231 = 11'he7 == fractionSum[12:2] ? 10'h12b : _GEN_230; // @[Multiplier.scala 64:55]
  assign _GEN_232 = 11'he8 == fractionSum[12:2] ? 10'h12c : _GEN_231; // @[Multiplier.scala 64:55]
  assign _GEN_233 = 11'he9 == fractionSum[12:2] ? 10'h12c : _GEN_232; // @[Multiplier.scala 64:55]
  assign _GEN_234 = 11'hea == fractionSum[12:2] ? 10'h12c : _GEN_233; // @[Multiplier.scala 64:55]
  assign _GEN_235 = 11'heb == fractionSum[12:2] ? 10'h12c : _GEN_234; // @[Multiplier.scala 64:55]
  assign _GEN_236 = 11'hec == fractionSum[12:2] ? 10'h12c : _GEN_235; // @[Multiplier.scala 64:55]
  assign _GEN_237 = 11'hed == fractionSum[12:2] ? 10'h12d : _GEN_236; // @[Multiplier.scala 64:55]
  assign _GEN_238 = 11'hee == fractionSum[12:2] ? 10'h12d : _GEN_237; // @[Multiplier.scala 64:55]
  assign _GEN_239 = 11'hef == fractionSum[12:2] ? 10'h12d : _GEN_238; // @[Multiplier.scala 64:55]
  assign _GEN_240 = 11'hf0 == fractionSum[12:2] ? 10'h12d : _GEN_239; // @[Multiplier.scala 64:55]
  assign _GEN_241 = 11'hf1 == fractionSum[12:2] ? 10'h12d : _GEN_240; // @[Multiplier.scala 64:55]
  assign _GEN_242 = 11'hf2 == fractionSum[12:2] ? 10'h12e : _GEN_241; // @[Multiplier.scala 64:55]
  assign _GEN_243 = 11'hf3 == fractionSum[12:2] ? 10'h12e : _GEN_242; // @[Multiplier.scala 64:55]
  assign _GEN_244 = 11'hf4 == fractionSum[12:2] ? 10'h12e : _GEN_243; // @[Multiplier.scala 64:55]
  assign _GEN_245 = 11'hf5 == fractionSum[12:2] ? 10'h12e : _GEN_244; // @[Multiplier.scala 64:55]
  assign _GEN_246 = 11'hf6 == fractionSum[12:2] ? 10'h12e : _GEN_245; // @[Multiplier.scala 64:55]
  assign _GEN_247 = 11'hf7 == fractionSum[12:2] ? 10'h12f : _GEN_246; // @[Multiplier.scala 64:55]
  assign _GEN_248 = 11'hf8 == fractionSum[12:2] ? 10'h12f : _GEN_247; // @[Multiplier.scala 64:55]
  assign _GEN_249 = 11'hf9 == fractionSum[12:2] ? 10'h12f : _GEN_248; // @[Multiplier.scala 64:55]
  assign _GEN_250 = 11'hfa == fractionSum[12:2] ? 10'h12f : _GEN_249; // @[Multiplier.scala 64:55]
  assign _GEN_251 = 11'hfb == fractionSum[12:2] ? 10'h12f : _GEN_250; // @[Multiplier.scala 64:55]
  assign _GEN_252 = 11'hfc == fractionSum[12:2] ? 10'h130 : _GEN_251; // @[Multiplier.scala 64:55]
  assign _GEN_253 = 11'hfd == fractionSum[12:2] ? 10'h130 : _GEN_252; // @[Multiplier.scala 64:55]
  assign _GEN_254 = 11'hfe == fractionSum[12:2] ? 10'h130 : _GEN_253; // @[Multiplier.scala 64:55]
  assign _GEN_255 = 11'hff == fractionSum[12:2] ? 10'h130 : _GEN_254; // @[Multiplier.scala 64:55]
  assign _GEN_256 = 11'h100 == fractionSum[12:2] ? 10'h130 : _GEN_255; // @[Multiplier.scala 64:55]
  assign _GEN_257 = 11'h101 == fractionSum[12:2] ? 10'h131 : _GEN_256; // @[Multiplier.scala 64:55]
  assign _GEN_258 = 11'h102 == fractionSum[12:2] ? 10'h131 : _GEN_257; // @[Multiplier.scala 64:55]
  assign _GEN_259 = 11'h103 == fractionSum[12:2] ? 10'h131 : _GEN_258; // @[Multiplier.scala 64:55]
  assign _GEN_260 = 11'h104 == fractionSum[12:2] ? 10'h131 : _GEN_259; // @[Multiplier.scala 64:55]
  assign _GEN_261 = 11'h105 == fractionSum[12:2] ? 10'h131 : _GEN_260; // @[Multiplier.scala 64:55]
  assign _GEN_262 = 11'h106 == fractionSum[12:2] ? 10'h132 : _GEN_261; // @[Multiplier.scala 64:55]
  assign _GEN_263 = 11'h107 == fractionSum[12:2] ? 10'h132 : _GEN_262; // @[Multiplier.scala 64:55]
  assign _GEN_264 = 11'h108 == fractionSum[12:2] ? 10'h132 : _GEN_263; // @[Multiplier.scala 64:55]
  assign _GEN_265 = 11'h109 == fractionSum[12:2] ? 10'h132 : _GEN_264; // @[Multiplier.scala 64:55]
  assign _GEN_266 = 11'h10a == fractionSum[12:2] ? 10'h133 : _GEN_265; // @[Multiplier.scala 64:55]
  assign _GEN_267 = 11'h10b == fractionSum[12:2] ? 10'h133 : _GEN_266; // @[Multiplier.scala 64:55]
  assign _GEN_268 = 11'h10c == fractionSum[12:2] ? 10'h133 : _GEN_267; // @[Multiplier.scala 64:55]
  assign _GEN_269 = 11'h10d == fractionSum[12:2] ? 10'h133 : _GEN_268; // @[Multiplier.scala 64:55]
  assign _GEN_270 = 11'h10e == fractionSum[12:2] ? 10'h133 : _GEN_269; // @[Multiplier.scala 64:55]
  assign _GEN_271 = 11'h10f == fractionSum[12:2] ? 10'h134 : _GEN_270; // @[Multiplier.scala 64:55]
  assign _GEN_272 = 11'h110 == fractionSum[12:2] ? 10'h134 : _GEN_271; // @[Multiplier.scala 64:55]
  assign _GEN_273 = 11'h111 == fractionSum[12:2] ? 10'h134 : _GEN_272; // @[Multiplier.scala 64:55]
  assign _GEN_274 = 11'h112 == fractionSum[12:2] ? 10'h134 : _GEN_273; // @[Multiplier.scala 64:55]
  assign _GEN_275 = 11'h113 == fractionSum[12:2] ? 10'h134 : _GEN_274; // @[Multiplier.scala 64:55]
  assign _GEN_276 = 11'h114 == fractionSum[12:2] ? 10'h135 : _GEN_275; // @[Multiplier.scala 64:55]
  assign _GEN_277 = 11'h115 == fractionSum[12:2] ? 10'h135 : _GEN_276; // @[Multiplier.scala 64:55]
  assign _GEN_278 = 11'h116 == fractionSum[12:2] ? 10'h135 : _GEN_277; // @[Multiplier.scala 64:55]
  assign _GEN_279 = 11'h117 == fractionSum[12:2] ? 10'h135 : _GEN_278; // @[Multiplier.scala 64:55]
  assign _GEN_280 = 11'h118 == fractionSum[12:2] ? 10'h135 : _GEN_279; // @[Multiplier.scala 64:55]
  assign _GEN_281 = 11'h119 == fractionSum[12:2] ? 10'h136 : _GEN_280; // @[Multiplier.scala 64:55]
  assign _GEN_282 = 11'h11a == fractionSum[12:2] ? 10'h136 : _GEN_281; // @[Multiplier.scala 64:55]
  assign _GEN_283 = 11'h11b == fractionSum[12:2] ? 10'h136 : _GEN_282; // @[Multiplier.scala 64:55]
  assign _GEN_284 = 11'h11c == fractionSum[12:2] ? 10'h136 : _GEN_283; // @[Multiplier.scala 64:55]
  assign _GEN_285 = 11'h11d == fractionSum[12:2] ? 10'h136 : _GEN_284; // @[Multiplier.scala 64:55]
  assign _GEN_286 = 11'h11e == fractionSum[12:2] ? 10'h137 : _GEN_285; // @[Multiplier.scala 64:55]
  assign _GEN_287 = 11'h11f == fractionSum[12:2] ? 10'h137 : _GEN_286; // @[Multiplier.scala 64:55]
  assign _GEN_288 = 11'h120 == fractionSum[12:2] ? 10'h137 : _GEN_287; // @[Multiplier.scala 64:55]
  assign _GEN_289 = 11'h121 == fractionSum[12:2] ? 10'h137 : _GEN_288; // @[Multiplier.scala 64:55]
  assign _GEN_290 = 11'h122 == fractionSum[12:2] ? 10'h138 : _GEN_289; // @[Multiplier.scala 64:55]
  assign _GEN_291 = 11'h123 == fractionSum[12:2] ? 10'h138 : _GEN_290; // @[Multiplier.scala 64:55]
  assign _GEN_292 = 11'h124 == fractionSum[12:2] ? 10'h138 : _GEN_291; // @[Multiplier.scala 64:55]
  assign _GEN_293 = 11'h125 == fractionSum[12:2] ? 10'h138 : _GEN_292; // @[Multiplier.scala 64:55]
  assign _GEN_294 = 11'h126 == fractionSum[12:2] ? 10'h138 : _GEN_293; // @[Multiplier.scala 64:55]
  assign _GEN_295 = 11'h127 == fractionSum[12:2] ? 10'h139 : _GEN_294; // @[Multiplier.scala 64:55]
  assign _GEN_296 = 11'h128 == fractionSum[12:2] ? 10'h139 : _GEN_295; // @[Multiplier.scala 64:55]
  assign _GEN_297 = 11'h129 == fractionSum[12:2] ? 10'h139 : _GEN_296; // @[Multiplier.scala 64:55]
  assign _GEN_298 = 11'h12a == fractionSum[12:2] ? 10'h139 : _GEN_297; // @[Multiplier.scala 64:55]
  assign _GEN_299 = 11'h12b == fractionSum[12:2] ? 10'h139 : _GEN_298; // @[Multiplier.scala 64:55]
  assign _GEN_300 = 11'h12c == fractionSum[12:2] ? 10'h13a : _GEN_299; // @[Multiplier.scala 64:55]
  assign _GEN_301 = 11'h12d == fractionSum[12:2] ? 10'h13a : _GEN_300; // @[Multiplier.scala 64:55]
  assign _GEN_302 = 11'h12e == fractionSum[12:2] ? 10'h13a : _GEN_301; // @[Multiplier.scala 64:55]
  assign _GEN_303 = 11'h12f == fractionSum[12:2] ? 10'h13a : _GEN_302; // @[Multiplier.scala 64:55]
  assign _GEN_304 = 11'h130 == fractionSum[12:2] ? 10'h13a : _GEN_303; // @[Multiplier.scala 64:55]
  assign _GEN_305 = 11'h131 == fractionSum[12:2] ? 10'h13b : _GEN_304; // @[Multiplier.scala 64:55]
  assign _GEN_306 = 11'h132 == fractionSum[12:2] ? 10'h13b : _GEN_305; // @[Multiplier.scala 64:55]
  assign _GEN_307 = 11'h133 == fractionSum[12:2] ? 10'h13b : _GEN_306; // @[Multiplier.scala 64:55]
  assign _GEN_308 = 11'h134 == fractionSum[12:2] ? 10'h13b : _GEN_307; // @[Multiplier.scala 64:55]
  assign _GEN_309 = 11'h135 == fractionSum[12:2] ? 10'h13c : _GEN_308; // @[Multiplier.scala 64:55]
  assign _GEN_310 = 11'h136 == fractionSum[12:2] ? 10'h13c : _GEN_309; // @[Multiplier.scala 64:55]
  assign _GEN_311 = 11'h137 == fractionSum[12:2] ? 10'h13c : _GEN_310; // @[Multiplier.scala 64:55]
  assign _GEN_312 = 11'h138 == fractionSum[12:2] ? 10'h13c : _GEN_311; // @[Multiplier.scala 64:55]
  assign _GEN_313 = 11'h139 == fractionSum[12:2] ? 10'h13c : _GEN_312; // @[Multiplier.scala 64:55]
  assign _GEN_314 = 11'h13a == fractionSum[12:2] ? 10'h13d : _GEN_313; // @[Multiplier.scala 64:55]
  assign _GEN_315 = 11'h13b == fractionSum[12:2] ? 10'h13d : _GEN_314; // @[Multiplier.scala 64:55]
  assign _GEN_316 = 11'h13c == fractionSum[12:2] ? 10'h13d : _GEN_315; // @[Multiplier.scala 64:55]
  assign _GEN_317 = 11'h13d == fractionSum[12:2] ? 10'h13d : _GEN_316; // @[Multiplier.scala 64:55]
  assign _GEN_318 = 11'h13e == fractionSum[12:2] ? 10'h13d : _GEN_317; // @[Multiplier.scala 64:55]
  assign _GEN_319 = 11'h13f == fractionSum[12:2] ? 10'h13e : _GEN_318; // @[Multiplier.scala 64:55]
  assign _GEN_320 = 11'h140 == fractionSum[12:2] ? 10'h13e : _GEN_319; // @[Multiplier.scala 64:55]
  assign _GEN_321 = 11'h141 == fractionSum[12:2] ? 10'h13e : _GEN_320; // @[Multiplier.scala 64:55]
  assign _GEN_322 = 11'h142 == fractionSum[12:2] ? 10'h13e : _GEN_321; // @[Multiplier.scala 64:55]
  assign _GEN_323 = 11'h143 == fractionSum[12:2] ? 10'h13f : _GEN_322; // @[Multiplier.scala 64:55]
  assign _GEN_324 = 11'h144 == fractionSum[12:2] ? 10'h13f : _GEN_323; // @[Multiplier.scala 64:55]
  assign _GEN_325 = 11'h145 == fractionSum[12:2] ? 10'h13f : _GEN_324; // @[Multiplier.scala 64:55]
  assign _GEN_326 = 11'h146 == fractionSum[12:2] ? 10'h13f : _GEN_325; // @[Multiplier.scala 64:55]
  assign _GEN_327 = 11'h147 == fractionSum[12:2] ? 10'h13f : _GEN_326; // @[Multiplier.scala 64:55]
  assign _GEN_328 = 11'h148 == fractionSum[12:2] ? 10'h140 : _GEN_327; // @[Multiplier.scala 64:55]
  assign _GEN_329 = 11'h149 == fractionSum[12:2] ? 10'h140 : _GEN_328; // @[Multiplier.scala 64:55]
  assign _GEN_330 = 11'h14a == fractionSum[12:2] ? 10'h140 : _GEN_329; // @[Multiplier.scala 64:55]
  assign _GEN_331 = 11'h14b == fractionSum[12:2] ? 10'h140 : _GEN_330; // @[Multiplier.scala 64:55]
  assign _GEN_332 = 11'h14c == fractionSum[12:2] ? 10'h141 : _GEN_331; // @[Multiplier.scala 64:55]
  assign _GEN_333 = 11'h14d == fractionSum[12:2] ? 10'h141 : _GEN_332; // @[Multiplier.scala 64:55]
  assign _GEN_334 = 11'h14e == fractionSum[12:2] ? 10'h141 : _GEN_333; // @[Multiplier.scala 64:55]
  assign _GEN_335 = 11'h14f == fractionSum[12:2] ? 10'h141 : _GEN_334; // @[Multiplier.scala 64:55]
  assign _GEN_336 = 11'h150 == fractionSum[12:2] ? 10'h141 : _GEN_335; // @[Multiplier.scala 64:55]
  assign _GEN_337 = 11'h151 == fractionSum[12:2] ? 10'h142 : _GEN_336; // @[Multiplier.scala 64:55]
  assign _GEN_338 = 11'h152 == fractionSum[12:2] ? 10'h142 : _GEN_337; // @[Multiplier.scala 64:55]
  assign _GEN_339 = 11'h153 == fractionSum[12:2] ? 10'h142 : _GEN_338; // @[Multiplier.scala 64:55]
  assign _GEN_340 = 11'h154 == fractionSum[12:2] ? 10'h142 : _GEN_339; // @[Multiplier.scala 64:55]
  assign _GEN_341 = 11'h155 == fractionSum[12:2] ? 10'h142 : _GEN_340; // @[Multiplier.scala 64:55]
  assign _GEN_342 = 11'h156 == fractionSum[12:2] ? 10'h143 : _GEN_341; // @[Multiplier.scala 64:55]
  assign _GEN_343 = 11'h157 == fractionSum[12:2] ? 10'h143 : _GEN_342; // @[Multiplier.scala 64:55]
  assign _GEN_344 = 11'h158 == fractionSum[12:2] ? 10'h143 : _GEN_343; // @[Multiplier.scala 64:55]
  assign _GEN_345 = 11'h159 == fractionSum[12:2] ? 10'h143 : _GEN_344; // @[Multiplier.scala 64:55]
  assign _GEN_346 = 11'h15a == fractionSum[12:2] ? 10'h144 : _GEN_345; // @[Multiplier.scala 64:55]
  assign _GEN_347 = 11'h15b == fractionSum[12:2] ? 10'h144 : _GEN_346; // @[Multiplier.scala 64:55]
  assign _GEN_348 = 11'h15c == fractionSum[12:2] ? 10'h144 : _GEN_347; // @[Multiplier.scala 64:55]
  assign _GEN_349 = 11'h15d == fractionSum[12:2] ? 10'h144 : _GEN_348; // @[Multiplier.scala 64:55]
  assign _GEN_350 = 11'h15e == fractionSum[12:2] ? 10'h144 : _GEN_349; // @[Multiplier.scala 64:55]
  assign _GEN_351 = 11'h15f == fractionSum[12:2] ? 10'h145 : _GEN_350; // @[Multiplier.scala 64:55]
  assign _GEN_352 = 11'h160 == fractionSum[12:2] ? 10'h145 : _GEN_351; // @[Multiplier.scala 64:55]
  assign _GEN_353 = 11'h161 == fractionSum[12:2] ? 10'h145 : _GEN_352; // @[Multiplier.scala 64:55]
  assign _GEN_354 = 11'h162 == fractionSum[12:2] ? 10'h145 : _GEN_353; // @[Multiplier.scala 64:55]
  assign _GEN_355 = 11'h163 == fractionSum[12:2] ? 10'h146 : _GEN_354; // @[Multiplier.scala 64:55]
  assign _GEN_356 = 11'h164 == fractionSum[12:2] ? 10'h146 : _GEN_355; // @[Multiplier.scala 64:55]
  assign _GEN_357 = 11'h165 == fractionSum[12:2] ? 10'h146 : _GEN_356; // @[Multiplier.scala 64:55]
  assign _GEN_358 = 11'h166 == fractionSum[12:2] ? 10'h146 : _GEN_357; // @[Multiplier.scala 64:55]
  assign _GEN_359 = 11'h167 == fractionSum[12:2] ? 10'h146 : _GEN_358; // @[Multiplier.scala 64:55]
  assign _GEN_360 = 11'h168 == fractionSum[12:2] ? 10'h147 : _GEN_359; // @[Multiplier.scala 64:55]
  assign _GEN_361 = 11'h169 == fractionSum[12:2] ? 10'h147 : _GEN_360; // @[Multiplier.scala 64:55]
  assign _GEN_362 = 11'h16a == fractionSum[12:2] ? 10'h147 : _GEN_361; // @[Multiplier.scala 64:55]
  assign _GEN_363 = 11'h16b == fractionSum[12:2] ? 10'h147 : _GEN_362; // @[Multiplier.scala 64:55]
  assign _GEN_364 = 11'h16c == fractionSum[12:2] ? 10'h148 : _GEN_363; // @[Multiplier.scala 64:55]
  assign _GEN_365 = 11'h16d == fractionSum[12:2] ? 10'h148 : _GEN_364; // @[Multiplier.scala 64:55]
  assign _GEN_366 = 11'h16e == fractionSum[12:2] ? 10'h148 : _GEN_365; // @[Multiplier.scala 64:55]
  assign _GEN_367 = 11'h16f == fractionSum[12:2] ? 10'h148 : _GEN_366; // @[Multiplier.scala 64:55]
  assign _GEN_368 = 11'h170 == fractionSum[12:2] ? 10'h148 : _GEN_367; // @[Multiplier.scala 64:55]
  assign _GEN_369 = 11'h171 == fractionSum[12:2] ? 10'h149 : _GEN_368; // @[Multiplier.scala 64:55]
  assign _GEN_370 = 11'h172 == fractionSum[12:2] ? 10'h149 : _GEN_369; // @[Multiplier.scala 64:55]
  assign _GEN_371 = 11'h173 == fractionSum[12:2] ? 10'h149 : _GEN_370; // @[Multiplier.scala 64:55]
  assign _GEN_372 = 11'h174 == fractionSum[12:2] ? 10'h149 : _GEN_371; // @[Multiplier.scala 64:55]
  assign _GEN_373 = 11'h175 == fractionSum[12:2] ? 10'h14a : _GEN_372; // @[Multiplier.scala 64:55]
  assign _GEN_374 = 11'h176 == fractionSum[12:2] ? 10'h14a : _GEN_373; // @[Multiplier.scala 64:55]
  assign _GEN_375 = 11'h177 == fractionSum[12:2] ? 10'h14a : _GEN_374; // @[Multiplier.scala 64:55]
  assign _GEN_376 = 11'h178 == fractionSum[12:2] ? 10'h14a : _GEN_375; // @[Multiplier.scala 64:55]
  assign _GEN_377 = 11'h179 == fractionSum[12:2] ? 10'h14a : _GEN_376; // @[Multiplier.scala 64:55]
  assign _GEN_378 = 11'h17a == fractionSum[12:2] ? 10'h14b : _GEN_377; // @[Multiplier.scala 64:55]
  assign _GEN_379 = 11'h17b == fractionSum[12:2] ? 10'h14b : _GEN_378; // @[Multiplier.scala 64:55]
  assign _GEN_380 = 11'h17c == fractionSum[12:2] ? 10'h14b : _GEN_379; // @[Multiplier.scala 64:55]
  assign _GEN_381 = 11'h17d == fractionSum[12:2] ? 10'h14b : _GEN_380; // @[Multiplier.scala 64:55]
  assign _GEN_382 = 11'h17e == fractionSum[12:2] ? 10'h14c : _GEN_381; // @[Multiplier.scala 64:55]
  assign _GEN_383 = 11'h17f == fractionSum[12:2] ? 10'h14c : _GEN_382; // @[Multiplier.scala 64:55]
  assign _GEN_384 = 11'h180 == fractionSum[12:2] ? 10'h14c : _GEN_383; // @[Multiplier.scala 64:55]
  assign _GEN_385 = 11'h181 == fractionSum[12:2] ? 10'h14c : _GEN_384; // @[Multiplier.scala 64:55]
  assign _GEN_386 = 11'h182 == fractionSum[12:2] ? 10'h14c : _GEN_385; // @[Multiplier.scala 64:55]
  assign _GEN_387 = 11'h183 == fractionSum[12:2] ? 10'h14d : _GEN_386; // @[Multiplier.scala 64:55]
  assign _GEN_388 = 11'h184 == fractionSum[12:2] ? 10'h14d : _GEN_387; // @[Multiplier.scala 64:55]
  assign _GEN_389 = 11'h185 == fractionSum[12:2] ? 10'h14d : _GEN_388; // @[Multiplier.scala 64:55]
  assign _GEN_390 = 11'h186 == fractionSum[12:2] ? 10'h14d : _GEN_389; // @[Multiplier.scala 64:55]
  assign _GEN_391 = 11'h187 == fractionSum[12:2] ? 10'h14e : _GEN_390; // @[Multiplier.scala 64:55]
  assign _GEN_392 = 11'h188 == fractionSum[12:2] ? 10'h14e : _GEN_391; // @[Multiplier.scala 64:55]
  assign _GEN_393 = 11'h189 == fractionSum[12:2] ? 10'h14e : _GEN_392; // @[Multiplier.scala 64:55]
  assign _GEN_394 = 11'h18a == fractionSum[12:2] ? 10'h14e : _GEN_393; // @[Multiplier.scala 64:55]
  assign _GEN_395 = 11'h18b == fractionSum[12:2] ? 10'h14e : _GEN_394; // @[Multiplier.scala 64:55]
  assign _GEN_396 = 11'h18c == fractionSum[12:2] ? 10'h14f : _GEN_395; // @[Multiplier.scala 64:55]
  assign _GEN_397 = 11'h18d == fractionSum[12:2] ? 10'h14f : _GEN_396; // @[Multiplier.scala 64:55]
  assign _GEN_398 = 11'h18e == fractionSum[12:2] ? 10'h14f : _GEN_397; // @[Multiplier.scala 64:55]
  assign _GEN_399 = 11'h18f == fractionSum[12:2] ? 10'h14f : _GEN_398; // @[Multiplier.scala 64:55]
  assign _GEN_400 = 11'h190 == fractionSum[12:2] ? 10'h150 : _GEN_399; // @[Multiplier.scala 64:55]
  assign _GEN_401 = 11'h191 == fractionSum[12:2] ? 10'h150 : _GEN_400; // @[Multiplier.scala 64:55]
  assign _GEN_402 = 11'h192 == fractionSum[12:2] ? 10'h150 : _GEN_401; // @[Multiplier.scala 64:55]
  assign _GEN_403 = 11'h193 == fractionSum[12:2] ? 10'h150 : _GEN_402; // @[Multiplier.scala 64:55]
  assign _GEN_404 = 11'h194 == fractionSum[12:2] ? 10'h151 : _GEN_403; // @[Multiplier.scala 64:55]
  assign _GEN_405 = 11'h195 == fractionSum[12:2] ? 10'h151 : _GEN_404; // @[Multiplier.scala 64:55]
  assign _GEN_406 = 11'h196 == fractionSum[12:2] ? 10'h151 : _GEN_405; // @[Multiplier.scala 64:55]
  assign _GEN_407 = 11'h197 == fractionSum[12:2] ? 10'h151 : _GEN_406; // @[Multiplier.scala 64:55]
  assign _GEN_408 = 11'h198 == fractionSum[12:2] ? 10'h151 : _GEN_407; // @[Multiplier.scala 64:55]
  assign _GEN_409 = 11'h199 == fractionSum[12:2] ? 10'h152 : _GEN_408; // @[Multiplier.scala 64:55]
  assign _GEN_410 = 11'h19a == fractionSum[12:2] ? 10'h152 : _GEN_409; // @[Multiplier.scala 64:55]
  assign _GEN_411 = 11'h19b == fractionSum[12:2] ? 10'h152 : _GEN_410; // @[Multiplier.scala 64:55]
  assign _GEN_412 = 11'h19c == fractionSum[12:2] ? 10'h152 : _GEN_411; // @[Multiplier.scala 64:55]
  assign _GEN_413 = 11'h19d == fractionSum[12:2] ? 10'h153 : _GEN_412; // @[Multiplier.scala 64:55]
  assign _GEN_414 = 11'h19e == fractionSum[12:2] ? 10'h153 : _GEN_413; // @[Multiplier.scala 64:55]
  assign _GEN_415 = 11'h19f == fractionSum[12:2] ? 10'h153 : _GEN_414; // @[Multiplier.scala 64:55]
  assign _GEN_416 = 11'h1a0 == fractionSum[12:2] ? 10'h153 : _GEN_415; // @[Multiplier.scala 64:55]
  assign _GEN_417 = 11'h1a1 == fractionSum[12:2] ? 10'h153 : _GEN_416; // @[Multiplier.scala 64:55]
  assign _GEN_418 = 11'h1a2 == fractionSum[12:2] ? 10'h154 : _GEN_417; // @[Multiplier.scala 64:55]
  assign _GEN_419 = 11'h1a3 == fractionSum[12:2] ? 10'h154 : _GEN_418; // @[Multiplier.scala 64:55]
  assign _GEN_420 = 11'h1a4 == fractionSum[12:2] ? 10'h154 : _GEN_419; // @[Multiplier.scala 64:55]
  assign _GEN_421 = 11'h1a5 == fractionSum[12:2] ? 10'h154 : _GEN_420; // @[Multiplier.scala 64:55]
  assign _GEN_422 = 11'h1a6 == fractionSum[12:2] ? 10'h155 : _GEN_421; // @[Multiplier.scala 64:55]
  assign _GEN_423 = 11'h1a7 == fractionSum[12:2] ? 10'h155 : _GEN_422; // @[Multiplier.scala 64:55]
  assign _GEN_424 = 11'h1a8 == fractionSum[12:2] ? 10'h155 : _GEN_423; // @[Multiplier.scala 64:55]
  assign _GEN_425 = 11'h1a9 == fractionSum[12:2] ? 10'h155 : _GEN_424; // @[Multiplier.scala 64:55]
  assign _GEN_426 = 11'h1aa == fractionSum[12:2] ? 10'h156 : _GEN_425; // @[Multiplier.scala 64:55]
  assign _GEN_427 = 11'h1ab == fractionSum[12:2] ? 10'h156 : _GEN_426; // @[Multiplier.scala 64:55]
  assign _GEN_428 = 11'h1ac == fractionSum[12:2] ? 10'h156 : _GEN_427; // @[Multiplier.scala 64:55]
  assign _GEN_429 = 11'h1ad == fractionSum[12:2] ? 10'h156 : _GEN_428; // @[Multiplier.scala 64:55]
  assign _GEN_430 = 11'h1ae == fractionSum[12:2] ? 10'h156 : _GEN_429; // @[Multiplier.scala 64:55]
  assign _GEN_431 = 11'h1af == fractionSum[12:2] ? 10'h157 : _GEN_430; // @[Multiplier.scala 64:55]
  assign _GEN_432 = 11'h1b0 == fractionSum[12:2] ? 10'h157 : _GEN_431; // @[Multiplier.scala 64:55]
  assign _GEN_433 = 11'h1b1 == fractionSum[12:2] ? 10'h157 : _GEN_432; // @[Multiplier.scala 64:55]
  assign _GEN_434 = 11'h1b2 == fractionSum[12:2] ? 10'h157 : _GEN_433; // @[Multiplier.scala 64:55]
  assign _GEN_435 = 11'h1b3 == fractionSum[12:2] ? 10'h158 : _GEN_434; // @[Multiplier.scala 64:55]
  assign _GEN_436 = 11'h1b4 == fractionSum[12:2] ? 10'h158 : _GEN_435; // @[Multiplier.scala 64:55]
  assign _GEN_437 = 11'h1b5 == fractionSum[12:2] ? 10'h158 : _GEN_436; // @[Multiplier.scala 64:55]
  assign _GEN_438 = 11'h1b6 == fractionSum[12:2] ? 10'h158 : _GEN_437; // @[Multiplier.scala 64:55]
  assign _GEN_439 = 11'h1b7 == fractionSum[12:2] ? 10'h159 : _GEN_438; // @[Multiplier.scala 64:55]
  assign _GEN_440 = 11'h1b8 == fractionSum[12:2] ? 10'h159 : _GEN_439; // @[Multiplier.scala 64:55]
  assign _GEN_441 = 11'h1b9 == fractionSum[12:2] ? 10'h159 : _GEN_440; // @[Multiplier.scala 64:55]
  assign _GEN_442 = 11'h1ba == fractionSum[12:2] ? 10'h159 : _GEN_441; // @[Multiplier.scala 64:55]
  assign _GEN_443 = 11'h1bb == fractionSum[12:2] ? 10'h15a : _GEN_442; // @[Multiplier.scala 64:55]
  assign _GEN_444 = 11'h1bc == fractionSum[12:2] ? 10'h15a : _GEN_443; // @[Multiplier.scala 64:55]
  assign _GEN_445 = 11'h1bd == fractionSum[12:2] ? 10'h15a : _GEN_444; // @[Multiplier.scala 64:55]
  assign _GEN_446 = 11'h1be == fractionSum[12:2] ? 10'h15a : _GEN_445; // @[Multiplier.scala 64:55]
  assign _GEN_447 = 11'h1bf == fractionSum[12:2] ? 10'h15a : _GEN_446; // @[Multiplier.scala 64:55]
  assign _GEN_448 = 11'h1c0 == fractionSum[12:2] ? 10'h15b : _GEN_447; // @[Multiplier.scala 64:55]
  assign _GEN_449 = 11'h1c1 == fractionSum[12:2] ? 10'h15b : _GEN_448; // @[Multiplier.scala 64:55]
  assign _GEN_450 = 11'h1c2 == fractionSum[12:2] ? 10'h15b : _GEN_449; // @[Multiplier.scala 64:55]
  assign _GEN_451 = 11'h1c3 == fractionSum[12:2] ? 10'h15b : _GEN_450; // @[Multiplier.scala 64:55]
  assign _GEN_452 = 11'h1c4 == fractionSum[12:2] ? 10'h15c : _GEN_451; // @[Multiplier.scala 64:55]
  assign _GEN_453 = 11'h1c5 == fractionSum[12:2] ? 10'h15c : _GEN_452; // @[Multiplier.scala 64:55]
  assign _GEN_454 = 11'h1c6 == fractionSum[12:2] ? 10'h15c : _GEN_453; // @[Multiplier.scala 64:55]
  assign _GEN_455 = 11'h1c7 == fractionSum[12:2] ? 10'h15c : _GEN_454; // @[Multiplier.scala 64:55]
  assign _GEN_456 = 11'h1c8 == fractionSum[12:2] ? 10'h15d : _GEN_455; // @[Multiplier.scala 64:55]
  assign _GEN_457 = 11'h1c9 == fractionSum[12:2] ? 10'h15d : _GEN_456; // @[Multiplier.scala 64:55]
  assign _GEN_458 = 11'h1ca == fractionSum[12:2] ? 10'h15d : _GEN_457; // @[Multiplier.scala 64:55]
  assign _GEN_459 = 11'h1cb == fractionSum[12:2] ? 10'h15d : _GEN_458; // @[Multiplier.scala 64:55]
  assign _GEN_460 = 11'h1cc == fractionSum[12:2] ? 10'h15e : _GEN_459; // @[Multiplier.scala 64:55]
  assign _GEN_461 = 11'h1cd == fractionSum[12:2] ? 10'h15e : _GEN_460; // @[Multiplier.scala 64:55]
  assign _GEN_462 = 11'h1ce == fractionSum[12:2] ? 10'h15e : _GEN_461; // @[Multiplier.scala 64:55]
  assign _GEN_463 = 11'h1cf == fractionSum[12:2] ? 10'h15e : _GEN_462; // @[Multiplier.scala 64:55]
  assign _GEN_464 = 11'h1d0 == fractionSum[12:2] ? 10'h15e : _GEN_463; // @[Multiplier.scala 64:55]
  assign _GEN_465 = 11'h1d1 == fractionSum[12:2] ? 10'h15f : _GEN_464; // @[Multiplier.scala 64:55]
  assign _GEN_466 = 11'h1d2 == fractionSum[12:2] ? 10'h15f : _GEN_465; // @[Multiplier.scala 64:55]
  assign _GEN_467 = 11'h1d3 == fractionSum[12:2] ? 10'h15f : _GEN_466; // @[Multiplier.scala 64:55]
  assign _GEN_468 = 11'h1d4 == fractionSum[12:2] ? 10'h15f : _GEN_467; // @[Multiplier.scala 64:55]
  assign _GEN_469 = 11'h1d5 == fractionSum[12:2] ? 10'h160 : _GEN_468; // @[Multiplier.scala 64:55]
  assign _GEN_470 = 11'h1d6 == fractionSum[12:2] ? 10'h160 : _GEN_469; // @[Multiplier.scala 64:55]
  assign _GEN_471 = 11'h1d7 == fractionSum[12:2] ? 10'h160 : _GEN_470; // @[Multiplier.scala 64:55]
  assign _GEN_472 = 11'h1d8 == fractionSum[12:2] ? 10'h160 : _GEN_471; // @[Multiplier.scala 64:55]
  assign _GEN_473 = 11'h1d9 == fractionSum[12:2] ? 10'h161 : _GEN_472; // @[Multiplier.scala 64:55]
  assign _GEN_474 = 11'h1da == fractionSum[12:2] ? 10'h161 : _GEN_473; // @[Multiplier.scala 64:55]
  assign _GEN_475 = 11'h1db == fractionSum[12:2] ? 10'h161 : _GEN_474; // @[Multiplier.scala 64:55]
  assign _GEN_476 = 11'h1dc == fractionSum[12:2] ? 10'h161 : _GEN_475; // @[Multiplier.scala 64:55]
  assign _GEN_477 = 11'h1dd == fractionSum[12:2] ? 10'h162 : _GEN_476; // @[Multiplier.scala 64:55]
  assign _GEN_478 = 11'h1de == fractionSum[12:2] ? 10'h162 : _GEN_477; // @[Multiplier.scala 64:55]
  assign _GEN_479 = 11'h1df == fractionSum[12:2] ? 10'h162 : _GEN_478; // @[Multiplier.scala 64:55]
  assign _GEN_480 = 11'h1e0 == fractionSum[12:2] ? 10'h162 : _GEN_479; // @[Multiplier.scala 64:55]
  assign _GEN_481 = 11'h1e1 == fractionSum[12:2] ? 10'h163 : _GEN_480; // @[Multiplier.scala 64:55]
  assign _GEN_482 = 11'h1e2 == fractionSum[12:2] ? 10'h163 : _GEN_481; // @[Multiplier.scala 64:55]
  assign _GEN_483 = 11'h1e3 == fractionSum[12:2] ? 10'h163 : _GEN_482; // @[Multiplier.scala 64:55]
  assign _GEN_484 = 11'h1e4 == fractionSum[12:2] ? 10'h163 : _GEN_483; // @[Multiplier.scala 64:55]
  assign _GEN_485 = 11'h1e5 == fractionSum[12:2] ? 10'h163 : _GEN_484; // @[Multiplier.scala 64:55]
  assign _GEN_486 = 11'h1e6 == fractionSum[12:2] ? 10'h164 : _GEN_485; // @[Multiplier.scala 64:55]
  assign _GEN_487 = 11'h1e7 == fractionSum[12:2] ? 10'h164 : _GEN_486; // @[Multiplier.scala 64:55]
  assign _GEN_488 = 11'h1e8 == fractionSum[12:2] ? 10'h164 : _GEN_487; // @[Multiplier.scala 64:55]
  assign _GEN_489 = 11'h1e9 == fractionSum[12:2] ? 10'h164 : _GEN_488; // @[Multiplier.scala 64:55]
  assign _GEN_490 = 11'h1ea == fractionSum[12:2] ? 10'h165 : _GEN_489; // @[Multiplier.scala 64:55]
  assign _GEN_491 = 11'h1eb == fractionSum[12:2] ? 10'h165 : _GEN_490; // @[Multiplier.scala 64:55]
  assign _GEN_492 = 11'h1ec == fractionSum[12:2] ? 10'h165 : _GEN_491; // @[Multiplier.scala 64:55]
  assign _GEN_493 = 11'h1ed == fractionSum[12:2] ? 10'h165 : _GEN_492; // @[Multiplier.scala 64:55]
  assign _GEN_494 = 11'h1ee == fractionSum[12:2] ? 10'h166 : _GEN_493; // @[Multiplier.scala 64:55]
  assign _GEN_495 = 11'h1ef == fractionSum[12:2] ? 10'h166 : _GEN_494; // @[Multiplier.scala 64:55]
  assign _GEN_496 = 11'h1f0 == fractionSum[12:2] ? 10'h166 : _GEN_495; // @[Multiplier.scala 64:55]
  assign _GEN_497 = 11'h1f1 == fractionSum[12:2] ? 10'h166 : _GEN_496; // @[Multiplier.scala 64:55]
  assign _GEN_498 = 11'h1f2 == fractionSum[12:2] ? 10'h167 : _GEN_497; // @[Multiplier.scala 64:55]
  assign _GEN_499 = 11'h1f3 == fractionSum[12:2] ? 10'h167 : _GEN_498; // @[Multiplier.scala 64:55]
  assign _GEN_500 = 11'h1f4 == fractionSum[12:2] ? 10'h167 : _GEN_499; // @[Multiplier.scala 64:55]
  assign _GEN_501 = 11'h1f5 == fractionSum[12:2] ? 10'h167 : _GEN_500; // @[Multiplier.scala 64:55]
  assign _GEN_502 = 11'h1f6 == fractionSum[12:2] ? 10'h168 : _GEN_501; // @[Multiplier.scala 64:55]
  assign _GEN_503 = 11'h1f7 == fractionSum[12:2] ? 10'h168 : _GEN_502; // @[Multiplier.scala 64:55]
  assign _GEN_504 = 11'h1f8 == fractionSum[12:2] ? 10'h168 : _GEN_503; // @[Multiplier.scala 64:55]
  assign _GEN_505 = 11'h1f9 == fractionSum[12:2] ? 10'h168 : _GEN_504; // @[Multiplier.scala 64:55]
  assign _GEN_506 = 11'h1fa == fractionSum[12:2] ? 10'h169 : _GEN_505; // @[Multiplier.scala 64:55]
  assign _GEN_507 = 11'h1fb == fractionSum[12:2] ? 10'h169 : _GEN_506; // @[Multiplier.scala 64:55]
  assign _GEN_508 = 11'h1fc == fractionSum[12:2] ? 10'h169 : _GEN_507; // @[Multiplier.scala 64:55]
  assign _GEN_509 = 11'h1fd == fractionSum[12:2] ? 10'h169 : _GEN_508; // @[Multiplier.scala 64:55]
  assign _GEN_510 = 11'h1fe == fractionSum[12:2] ? 10'h16a : _GEN_509; // @[Multiplier.scala 64:55]
  assign _GEN_511 = 11'h1ff == fractionSum[12:2] ? 10'h16a : _GEN_510; // @[Multiplier.scala 64:55]
  assign _GEN_512 = 11'h200 == fractionSum[12:2] ? 10'h16a : _GEN_511; // @[Multiplier.scala 64:55]
  assign _GEN_513 = 11'h201 == fractionSum[12:2] ? 10'h16a : _GEN_512; // @[Multiplier.scala 64:55]
  assign _GEN_514 = 11'h202 == fractionSum[12:2] ? 10'h16b : _GEN_513; // @[Multiplier.scala 64:55]
  assign _GEN_515 = 11'h203 == fractionSum[12:2] ? 10'h16b : _GEN_514; // @[Multiplier.scala 64:55]
  assign _GEN_516 = 11'h204 == fractionSum[12:2] ? 10'h16b : _GEN_515; // @[Multiplier.scala 64:55]
  assign _GEN_517 = 11'h205 == fractionSum[12:2] ? 10'h16b : _GEN_516; // @[Multiplier.scala 64:55]
  assign _GEN_518 = 11'h206 == fractionSum[12:2] ? 10'h16c : _GEN_517; // @[Multiplier.scala 64:55]
  assign _GEN_519 = 11'h207 == fractionSum[12:2] ? 10'h16c : _GEN_518; // @[Multiplier.scala 64:55]
  assign _GEN_520 = 11'h208 == fractionSum[12:2] ? 10'h16c : _GEN_519; // @[Multiplier.scala 64:55]
  assign _GEN_521 = 11'h209 == fractionSum[12:2] ? 10'h16c : _GEN_520; // @[Multiplier.scala 64:55]
  assign _GEN_522 = 11'h20a == fractionSum[12:2] ? 10'h16c : _GEN_521; // @[Multiplier.scala 64:55]
  assign _GEN_523 = 11'h20b == fractionSum[12:2] ? 10'h16d : _GEN_522; // @[Multiplier.scala 64:55]
  assign _GEN_524 = 11'h20c == fractionSum[12:2] ? 10'h16d : _GEN_523; // @[Multiplier.scala 64:55]
  assign _GEN_525 = 11'h20d == fractionSum[12:2] ? 10'h16d : _GEN_524; // @[Multiplier.scala 64:55]
  assign _GEN_526 = 11'h20e == fractionSum[12:2] ? 10'h16d : _GEN_525; // @[Multiplier.scala 64:55]
  assign _GEN_527 = 11'h20f == fractionSum[12:2] ? 10'h16e : _GEN_526; // @[Multiplier.scala 64:55]
  assign _GEN_528 = 11'h210 == fractionSum[12:2] ? 10'h16e : _GEN_527; // @[Multiplier.scala 64:55]
  assign _GEN_529 = 11'h211 == fractionSum[12:2] ? 10'h16e : _GEN_528; // @[Multiplier.scala 64:55]
  assign _GEN_530 = 11'h212 == fractionSum[12:2] ? 10'h16e : _GEN_529; // @[Multiplier.scala 64:55]
  assign _GEN_531 = 11'h213 == fractionSum[12:2] ? 10'h16f : _GEN_530; // @[Multiplier.scala 64:55]
  assign _GEN_532 = 11'h214 == fractionSum[12:2] ? 10'h16f : _GEN_531; // @[Multiplier.scala 64:55]
  assign _GEN_533 = 11'h215 == fractionSum[12:2] ? 10'h16f : _GEN_532; // @[Multiplier.scala 64:55]
  assign _GEN_534 = 11'h216 == fractionSum[12:2] ? 10'h16f : _GEN_533; // @[Multiplier.scala 64:55]
  assign _GEN_535 = 11'h217 == fractionSum[12:2] ? 10'h170 : _GEN_534; // @[Multiplier.scala 64:55]
  assign _GEN_536 = 11'h218 == fractionSum[12:2] ? 10'h170 : _GEN_535; // @[Multiplier.scala 64:55]
  assign _GEN_537 = 11'h219 == fractionSum[12:2] ? 10'h170 : _GEN_536; // @[Multiplier.scala 64:55]
  assign _GEN_538 = 11'h21a == fractionSum[12:2] ? 10'h170 : _GEN_537; // @[Multiplier.scala 64:55]
  assign _GEN_539 = 11'h21b == fractionSum[12:2] ? 10'h171 : _GEN_538; // @[Multiplier.scala 64:55]
  assign _GEN_540 = 11'h21c == fractionSum[12:2] ? 10'h171 : _GEN_539; // @[Multiplier.scala 64:55]
  assign _GEN_541 = 11'h21d == fractionSum[12:2] ? 10'h171 : _GEN_540; // @[Multiplier.scala 64:55]
  assign _GEN_542 = 11'h21e == fractionSum[12:2] ? 10'h171 : _GEN_541; // @[Multiplier.scala 64:55]
  assign _GEN_543 = 11'h21f == fractionSum[12:2] ? 10'h172 : _GEN_542; // @[Multiplier.scala 64:55]
  assign _GEN_544 = 11'h220 == fractionSum[12:2] ? 10'h172 : _GEN_543; // @[Multiplier.scala 64:55]
  assign _GEN_545 = 11'h221 == fractionSum[12:2] ? 10'h172 : _GEN_544; // @[Multiplier.scala 64:55]
  assign _GEN_546 = 11'h222 == fractionSum[12:2] ? 10'h172 : _GEN_545; // @[Multiplier.scala 64:55]
  assign _GEN_547 = 11'h223 == fractionSum[12:2] ? 10'h173 : _GEN_546; // @[Multiplier.scala 64:55]
  assign _GEN_548 = 11'h224 == fractionSum[12:2] ? 10'h173 : _GEN_547; // @[Multiplier.scala 64:55]
  assign _GEN_549 = 11'h225 == fractionSum[12:2] ? 10'h173 : _GEN_548; // @[Multiplier.scala 64:55]
  assign _GEN_550 = 11'h226 == fractionSum[12:2] ? 10'h173 : _GEN_549; // @[Multiplier.scala 64:55]
  assign _GEN_551 = 11'h227 == fractionSum[12:2] ? 10'h174 : _GEN_550; // @[Multiplier.scala 64:55]
  assign _GEN_552 = 11'h228 == fractionSum[12:2] ? 10'h174 : _GEN_551; // @[Multiplier.scala 64:55]
  assign _GEN_553 = 11'h229 == fractionSum[12:2] ? 10'h174 : _GEN_552; // @[Multiplier.scala 64:55]
  assign _GEN_554 = 11'h22a == fractionSum[12:2] ? 10'h174 : _GEN_553; // @[Multiplier.scala 64:55]
  assign _GEN_555 = 11'h22b == fractionSum[12:2] ? 10'h175 : _GEN_554; // @[Multiplier.scala 64:55]
  assign _GEN_556 = 11'h22c == fractionSum[12:2] ? 10'h175 : _GEN_555; // @[Multiplier.scala 64:55]
  assign _GEN_557 = 11'h22d == fractionSum[12:2] ? 10'h175 : _GEN_556; // @[Multiplier.scala 64:55]
  assign _GEN_558 = 11'h22e == fractionSum[12:2] ? 10'h175 : _GEN_557; // @[Multiplier.scala 64:55]
  assign _GEN_559 = 11'h22f == fractionSum[12:2] ? 10'h176 : _GEN_558; // @[Multiplier.scala 64:55]
  assign _GEN_560 = 11'h230 == fractionSum[12:2] ? 10'h176 : _GEN_559; // @[Multiplier.scala 64:55]
  assign _GEN_561 = 11'h231 == fractionSum[12:2] ? 10'h176 : _GEN_560; // @[Multiplier.scala 64:55]
  assign _GEN_562 = 11'h232 == fractionSum[12:2] ? 10'h177 : _GEN_561; // @[Multiplier.scala 64:55]
  assign _GEN_563 = 11'h233 == fractionSum[12:2] ? 10'h177 : _GEN_562; // @[Multiplier.scala 64:55]
  assign _GEN_564 = 11'h234 == fractionSum[12:2] ? 10'h177 : _GEN_563; // @[Multiplier.scala 64:55]
  assign _GEN_565 = 11'h235 == fractionSum[12:2] ? 10'h177 : _GEN_564; // @[Multiplier.scala 64:55]
  assign _GEN_566 = 11'h236 == fractionSum[12:2] ? 10'h178 : _GEN_565; // @[Multiplier.scala 64:55]
  assign _GEN_567 = 11'h237 == fractionSum[12:2] ? 10'h178 : _GEN_566; // @[Multiplier.scala 64:55]
  assign _GEN_568 = 11'h238 == fractionSum[12:2] ? 10'h178 : _GEN_567; // @[Multiplier.scala 64:55]
  assign _GEN_569 = 11'h239 == fractionSum[12:2] ? 10'h178 : _GEN_568; // @[Multiplier.scala 64:55]
  assign _GEN_570 = 11'h23a == fractionSum[12:2] ? 10'h179 : _GEN_569; // @[Multiplier.scala 64:55]
  assign _GEN_571 = 11'h23b == fractionSum[12:2] ? 10'h179 : _GEN_570; // @[Multiplier.scala 64:55]
  assign _GEN_572 = 11'h23c == fractionSum[12:2] ? 10'h179 : _GEN_571; // @[Multiplier.scala 64:55]
  assign _GEN_573 = 11'h23d == fractionSum[12:2] ? 10'h179 : _GEN_572; // @[Multiplier.scala 64:55]
  assign _GEN_574 = 11'h23e == fractionSum[12:2] ? 10'h17a : _GEN_573; // @[Multiplier.scala 64:55]
  assign _GEN_575 = 11'h23f == fractionSum[12:2] ? 10'h17a : _GEN_574; // @[Multiplier.scala 64:55]
  assign _GEN_576 = 11'h240 == fractionSum[12:2] ? 10'h17a : _GEN_575; // @[Multiplier.scala 64:55]
  assign _GEN_577 = 11'h241 == fractionSum[12:2] ? 10'h17a : _GEN_576; // @[Multiplier.scala 64:55]
  assign _GEN_578 = 11'h242 == fractionSum[12:2] ? 10'h17b : _GEN_577; // @[Multiplier.scala 64:55]
  assign _GEN_579 = 11'h243 == fractionSum[12:2] ? 10'h17b : _GEN_578; // @[Multiplier.scala 64:55]
  assign _GEN_580 = 11'h244 == fractionSum[12:2] ? 10'h17b : _GEN_579; // @[Multiplier.scala 64:55]
  assign _GEN_581 = 11'h245 == fractionSum[12:2] ? 10'h17b : _GEN_580; // @[Multiplier.scala 64:55]
  assign _GEN_582 = 11'h246 == fractionSum[12:2] ? 10'h17c : _GEN_581; // @[Multiplier.scala 64:55]
  assign _GEN_583 = 11'h247 == fractionSum[12:2] ? 10'h17c : _GEN_582; // @[Multiplier.scala 64:55]
  assign _GEN_584 = 11'h248 == fractionSum[12:2] ? 10'h17c : _GEN_583; // @[Multiplier.scala 64:55]
  assign _GEN_585 = 11'h249 == fractionSum[12:2] ? 10'h17c : _GEN_584; // @[Multiplier.scala 64:55]
  assign _GEN_586 = 11'h24a == fractionSum[12:2] ? 10'h17d : _GEN_585; // @[Multiplier.scala 64:55]
  assign _GEN_587 = 11'h24b == fractionSum[12:2] ? 10'h17d : _GEN_586; // @[Multiplier.scala 64:55]
  assign _GEN_588 = 11'h24c == fractionSum[12:2] ? 10'h17d : _GEN_587; // @[Multiplier.scala 64:55]
  assign _GEN_589 = 11'h24d == fractionSum[12:2] ? 10'h17d : _GEN_588; // @[Multiplier.scala 64:55]
  assign _GEN_590 = 11'h24e == fractionSum[12:2] ? 10'h17e : _GEN_589; // @[Multiplier.scala 64:55]
  assign _GEN_591 = 11'h24f == fractionSum[12:2] ? 10'h17e : _GEN_590; // @[Multiplier.scala 64:55]
  assign _GEN_592 = 11'h250 == fractionSum[12:2] ? 10'h17e : _GEN_591; // @[Multiplier.scala 64:55]
  assign _GEN_593 = 11'h251 == fractionSum[12:2] ? 10'h17e : _GEN_592; // @[Multiplier.scala 64:55]
  assign _GEN_594 = 11'h252 == fractionSum[12:2] ? 10'h17f : _GEN_593; // @[Multiplier.scala 64:55]
  assign _GEN_595 = 11'h253 == fractionSum[12:2] ? 10'h17f : _GEN_594; // @[Multiplier.scala 64:55]
  assign _GEN_596 = 11'h254 == fractionSum[12:2] ? 10'h17f : _GEN_595; // @[Multiplier.scala 64:55]
  assign _GEN_597 = 11'h255 == fractionSum[12:2] ? 10'h17f : _GEN_596; // @[Multiplier.scala 64:55]
  assign _GEN_598 = 11'h256 == fractionSum[12:2] ? 10'h180 : _GEN_597; // @[Multiplier.scala 64:55]
  assign _GEN_599 = 11'h257 == fractionSum[12:2] ? 10'h180 : _GEN_598; // @[Multiplier.scala 64:55]
  assign _GEN_600 = 11'h258 == fractionSum[12:2] ? 10'h180 : _GEN_599; // @[Multiplier.scala 64:55]
  assign _GEN_601 = 11'h259 == fractionSum[12:2] ? 10'h181 : _GEN_600; // @[Multiplier.scala 64:55]
  assign _GEN_602 = 11'h25a == fractionSum[12:2] ? 10'h181 : _GEN_601; // @[Multiplier.scala 64:55]
  assign _GEN_603 = 11'h25b == fractionSum[12:2] ? 10'h181 : _GEN_602; // @[Multiplier.scala 64:55]
  assign _GEN_604 = 11'h25c == fractionSum[12:2] ? 10'h181 : _GEN_603; // @[Multiplier.scala 64:55]
  assign _GEN_605 = 11'h25d == fractionSum[12:2] ? 10'h182 : _GEN_604; // @[Multiplier.scala 64:55]
  assign _GEN_606 = 11'h25e == fractionSum[12:2] ? 10'h182 : _GEN_605; // @[Multiplier.scala 64:55]
  assign _GEN_607 = 11'h25f == fractionSum[12:2] ? 10'h182 : _GEN_606; // @[Multiplier.scala 64:55]
  assign _GEN_608 = 11'h260 == fractionSum[12:2] ? 10'h182 : _GEN_607; // @[Multiplier.scala 64:55]
  assign _GEN_609 = 11'h261 == fractionSum[12:2] ? 10'h183 : _GEN_608; // @[Multiplier.scala 64:55]
  assign _GEN_610 = 11'h262 == fractionSum[12:2] ? 10'h183 : _GEN_609; // @[Multiplier.scala 64:55]
  assign _GEN_611 = 11'h263 == fractionSum[12:2] ? 10'h183 : _GEN_610; // @[Multiplier.scala 64:55]
  assign _GEN_612 = 11'h264 == fractionSum[12:2] ? 10'h183 : _GEN_611; // @[Multiplier.scala 64:55]
  assign _GEN_613 = 11'h265 == fractionSum[12:2] ? 10'h184 : _GEN_612; // @[Multiplier.scala 64:55]
  assign _GEN_614 = 11'h266 == fractionSum[12:2] ? 10'h184 : _GEN_613; // @[Multiplier.scala 64:55]
  assign _GEN_615 = 11'h267 == fractionSum[12:2] ? 10'h184 : _GEN_614; // @[Multiplier.scala 64:55]
  assign _GEN_616 = 11'h268 == fractionSum[12:2] ? 10'h184 : _GEN_615; // @[Multiplier.scala 64:55]
  assign _GEN_617 = 11'h269 == fractionSum[12:2] ? 10'h185 : _GEN_616; // @[Multiplier.scala 64:55]
  assign _GEN_618 = 11'h26a == fractionSum[12:2] ? 10'h185 : _GEN_617; // @[Multiplier.scala 64:55]
  assign _GEN_619 = 11'h26b == fractionSum[12:2] ? 10'h185 : _GEN_618; // @[Multiplier.scala 64:55]
  assign _GEN_620 = 11'h26c == fractionSum[12:2] ? 10'h185 : _GEN_619; // @[Multiplier.scala 64:55]
  assign _GEN_621 = 11'h26d == fractionSum[12:2] ? 10'h186 : _GEN_620; // @[Multiplier.scala 64:55]
  assign _GEN_622 = 11'h26e == fractionSum[12:2] ? 10'h186 : _GEN_621; // @[Multiplier.scala 64:55]
  assign _GEN_623 = 11'h26f == fractionSum[12:2] ? 10'h186 : _GEN_622; // @[Multiplier.scala 64:55]
  assign _GEN_624 = 11'h270 == fractionSum[12:2] ? 10'h187 : _GEN_623; // @[Multiplier.scala 64:55]
  assign _GEN_625 = 11'h271 == fractionSum[12:2] ? 10'h187 : _GEN_624; // @[Multiplier.scala 64:55]
  assign _GEN_626 = 11'h272 == fractionSum[12:2] ? 10'h187 : _GEN_625; // @[Multiplier.scala 64:55]
  assign _GEN_627 = 11'h273 == fractionSum[12:2] ? 10'h187 : _GEN_626; // @[Multiplier.scala 64:55]
  assign _GEN_628 = 11'h274 == fractionSum[12:2] ? 10'h188 : _GEN_627; // @[Multiplier.scala 64:55]
  assign _GEN_629 = 11'h275 == fractionSum[12:2] ? 10'h188 : _GEN_628; // @[Multiplier.scala 64:55]
  assign _GEN_630 = 11'h276 == fractionSum[12:2] ? 10'h188 : _GEN_629; // @[Multiplier.scala 64:55]
  assign _GEN_631 = 11'h277 == fractionSum[12:2] ? 10'h188 : _GEN_630; // @[Multiplier.scala 64:55]
  assign _GEN_632 = 11'h278 == fractionSum[12:2] ? 10'h189 : _GEN_631; // @[Multiplier.scala 64:55]
  assign _GEN_633 = 11'h279 == fractionSum[12:2] ? 10'h189 : _GEN_632; // @[Multiplier.scala 64:55]
  assign _GEN_634 = 11'h27a == fractionSum[12:2] ? 10'h189 : _GEN_633; // @[Multiplier.scala 64:55]
  assign _GEN_635 = 11'h27b == fractionSum[12:2] ? 10'h189 : _GEN_634; // @[Multiplier.scala 64:55]
  assign _GEN_636 = 11'h27c == fractionSum[12:2] ? 10'h18a : _GEN_635; // @[Multiplier.scala 64:55]
  assign _GEN_637 = 11'h27d == fractionSum[12:2] ? 10'h18a : _GEN_636; // @[Multiplier.scala 64:55]
  assign _GEN_638 = 11'h27e == fractionSum[12:2] ? 10'h18a : _GEN_637; // @[Multiplier.scala 64:55]
  assign _GEN_639 = 11'h27f == fractionSum[12:2] ? 10'h18b : _GEN_638; // @[Multiplier.scala 64:55]
  assign _GEN_640 = 11'h280 == fractionSum[12:2] ? 10'h18b : _GEN_639; // @[Multiplier.scala 64:55]
  assign _GEN_641 = 11'h281 == fractionSum[12:2] ? 10'h18b : _GEN_640; // @[Multiplier.scala 64:55]
  assign _GEN_642 = 11'h282 == fractionSum[12:2] ? 10'h18b : _GEN_641; // @[Multiplier.scala 64:55]
  assign _GEN_643 = 11'h283 == fractionSum[12:2] ? 10'h18c : _GEN_642; // @[Multiplier.scala 64:55]
  assign _GEN_644 = 11'h284 == fractionSum[12:2] ? 10'h18c : _GEN_643; // @[Multiplier.scala 64:55]
  assign _GEN_645 = 11'h285 == fractionSum[12:2] ? 10'h18c : _GEN_644; // @[Multiplier.scala 64:55]
  assign _GEN_646 = 11'h286 == fractionSum[12:2] ? 10'h18c : _GEN_645; // @[Multiplier.scala 64:55]
  assign _GEN_647 = 11'h287 == fractionSum[12:2] ? 10'h18d : _GEN_646; // @[Multiplier.scala 64:55]
  assign _GEN_648 = 11'h288 == fractionSum[12:2] ? 10'h18d : _GEN_647; // @[Multiplier.scala 64:55]
  assign _GEN_649 = 11'h289 == fractionSum[12:2] ? 10'h18d : _GEN_648; // @[Multiplier.scala 64:55]
  assign _GEN_650 = 11'h28a == fractionSum[12:2] ? 10'h18d : _GEN_649; // @[Multiplier.scala 64:55]
  assign _GEN_651 = 11'h28b == fractionSum[12:2] ? 10'h18e : _GEN_650; // @[Multiplier.scala 64:55]
  assign _GEN_652 = 11'h28c == fractionSum[12:2] ? 10'h18e : _GEN_651; // @[Multiplier.scala 64:55]
  assign _GEN_653 = 11'h28d == fractionSum[12:2] ? 10'h18e : _GEN_652; // @[Multiplier.scala 64:55]
  assign _GEN_654 = 11'h28e == fractionSum[12:2] ? 10'h18f : _GEN_653; // @[Multiplier.scala 64:55]
  assign _GEN_655 = 11'h28f == fractionSum[12:2] ? 10'h18f : _GEN_654; // @[Multiplier.scala 64:55]
  assign _GEN_656 = 11'h290 == fractionSum[12:2] ? 10'h18f : _GEN_655; // @[Multiplier.scala 64:55]
  assign _GEN_657 = 11'h291 == fractionSum[12:2] ? 10'h18f : _GEN_656; // @[Multiplier.scala 64:55]
  assign _GEN_658 = 11'h292 == fractionSum[12:2] ? 10'h190 : _GEN_657; // @[Multiplier.scala 64:55]
  assign _GEN_659 = 11'h293 == fractionSum[12:2] ? 10'h190 : _GEN_658; // @[Multiplier.scala 64:55]
  assign _GEN_660 = 11'h294 == fractionSum[12:2] ? 10'h190 : _GEN_659; // @[Multiplier.scala 64:55]
  assign _GEN_661 = 11'h295 == fractionSum[12:2] ? 10'h190 : _GEN_660; // @[Multiplier.scala 64:55]
  assign _GEN_662 = 11'h296 == fractionSum[12:2] ? 10'h191 : _GEN_661; // @[Multiplier.scala 64:55]
  assign _GEN_663 = 11'h297 == fractionSum[12:2] ? 10'h191 : _GEN_662; // @[Multiplier.scala 64:55]
  assign _GEN_664 = 11'h298 == fractionSum[12:2] ? 10'h191 : _GEN_663; // @[Multiplier.scala 64:55]
  assign _GEN_665 = 11'h299 == fractionSum[12:2] ? 10'h192 : _GEN_664; // @[Multiplier.scala 64:55]
  assign _GEN_666 = 11'h29a == fractionSum[12:2] ? 10'h192 : _GEN_665; // @[Multiplier.scala 64:55]
  assign _GEN_667 = 11'h29b == fractionSum[12:2] ? 10'h192 : _GEN_666; // @[Multiplier.scala 64:55]
  assign _GEN_668 = 11'h29c == fractionSum[12:2] ? 10'h192 : _GEN_667; // @[Multiplier.scala 64:55]
  assign _GEN_669 = 11'h29d == fractionSum[12:2] ? 10'h193 : _GEN_668; // @[Multiplier.scala 64:55]
  assign _GEN_670 = 11'h29e == fractionSum[12:2] ? 10'h193 : _GEN_669; // @[Multiplier.scala 64:55]
  assign _GEN_671 = 11'h29f == fractionSum[12:2] ? 10'h193 : _GEN_670; // @[Multiplier.scala 64:55]
  assign _GEN_672 = 11'h2a0 == fractionSum[12:2] ? 10'h193 : _GEN_671; // @[Multiplier.scala 64:55]
  assign _GEN_673 = 11'h2a1 == fractionSum[12:2] ? 10'h194 : _GEN_672; // @[Multiplier.scala 64:55]
  assign _GEN_674 = 11'h2a2 == fractionSum[12:2] ? 10'h194 : _GEN_673; // @[Multiplier.scala 64:55]
  assign _GEN_675 = 11'h2a3 == fractionSum[12:2] ? 10'h194 : _GEN_674; // @[Multiplier.scala 64:55]
  assign _GEN_676 = 11'h2a4 == fractionSum[12:2] ? 10'h195 : _GEN_675; // @[Multiplier.scala 64:55]
  assign _GEN_677 = 11'h2a5 == fractionSum[12:2] ? 10'h195 : _GEN_676; // @[Multiplier.scala 64:55]
  assign _GEN_678 = 11'h2a6 == fractionSum[12:2] ? 10'h195 : _GEN_677; // @[Multiplier.scala 64:55]
  assign _GEN_679 = 11'h2a7 == fractionSum[12:2] ? 10'h195 : _GEN_678; // @[Multiplier.scala 64:55]
  assign _GEN_680 = 11'h2a8 == fractionSum[12:2] ? 10'h196 : _GEN_679; // @[Multiplier.scala 64:55]
  assign _GEN_681 = 11'h2a9 == fractionSum[12:2] ? 10'h196 : _GEN_680; // @[Multiplier.scala 64:55]
  assign _GEN_682 = 11'h2aa == fractionSum[12:2] ? 10'h196 : _GEN_681; // @[Multiplier.scala 64:55]
  assign _GEN_683 = 11'h2ab == fractionSum[12:2] ? 10'h196 : _GEN_682; // @[Multiplier.scala 64:55]
  assign _GEN_684 = 11'h2ac == fractionSum[12:2] ? 10'h197 : _GEN_683; // @[Multiplier.scala 64:55]
  assign _GEN_685 = 11'h2ad == fractionSum[12:2] ? 10'h197 : _GEN_684; // @[Multiplier.scala 64:55]
  assign _GEN_686 = 11'h2ae == fractionSum[12:2] ? 10'h197 : _GEN_685; // @[Multiplier.scala 64:55]
  assign _GEN_687 = 11'h2af == fractionSum[12:2] ? 10'h198 : _GEN_686; // @[Multiplier.scala 64:55]
  assign _GEN_688 = 11'h2b0 == fractionSum[12:2] ? 10'h198 : _GEN_687; // @[Multiplier.scala 64:55]
  assign _GEN_689 = 11'h2b1 == fractionSum[12:2] ? 10'h198 : _GEN_688; // @[Multiplier.scala 64:55]
  assign _GEN_690 = 11'h2b2 == fractionSum[12:2] ? 10'h198 : _GEN_689; // @[Multiplier.scala 64:55]
  assign _GEN_691 = 11'h2b3 == fractionSum[12:2] ? 10'h199 : _GEN_690; // @[Multiplier.scala 64:55]
  assign _GEN_692 = 11'h2b4 == fractionSum[12:2] ? 10'h199 : _GEN_691; // @[Multiplier.scala 64:55]
  assign _GEN_693 = 11'h2b5 == fractionSum[12:2] ? 10'h199 : _GEN_692; // @[Multiplier.scala 64:55]
  assign _GEN_694 = 11'h2b6 == fractionSum[12:2] ? 10'h19a : _GEN_693; // @[Multiplier.scala 64:55]
  assign _GEN_695 = 11'h2b7 == fractionSum[12:2] ? 10'h19a : _GEN_694; // @[Multiplier.scala 64:55]
  assign _GEN_696 = 11'h2b8 == fractionSum[12:2] ? 10'h19a : _GEN_695; // @[Multiplier.scala 64:55]
  assign _GEN_697 = 11'h2b9 == fractionSum[12:2] ? 10'h19a : _GEN_696; // @[Multiplier.scala 64:55]
  assign _GEN_698 = 11'h2ba == fractionSum[12:2] ? 10'h19b : _GEN_697; // @[Multiplier.scala 64:55]
  assign _GEN_699 = 11'h2bb == fractionSum[12:2] ? 10'h19b : _GEN_698; // @[Multiplier.scala 64:55]
  assign _GEN_700 = 11'h2bc == fractionSum[12:2] ? 10'h19b : _GEN_699; // @[Multiplier.scala 64:55]
  assign _GEN_701 = 11'h2bd == fractionSum[12:2] ? 10'h19b : _GEN_700; // @[Multiplier.scala 64:55]
  assign _GEN_702 = 11'h2be == fractionSum[12:2] ? 10'h19c : _GEN_701; // @[Multiplier.scala 64:55]
  assign _GEN_703 = 11'h2bf == fractionSum[12:2] ? 10'h19c : _GEN_702; // @[Multiplier.scala 64:55]
  assign _GEN_704 = 11'h2c0 == fractionSum[12:2] ? 10'h19c : _GEN_703; // @[Multiplier.scala 64:55]
  assign _GEN_705 = 11'h2c1 == fractionSum[12:2] ? 10'h19d : _GEN_704; // @[Multiplier.scala 64:55]
  assign _GEN_706 = 11'h2c2 == fractionSum[12:2] ? 10'h19d : _GEN_705; // @[Multiplier.scala 64:55]
  assign _GEN_707 = 11'h2c3 == fractionSum[12:2] ? 10'h19d : _GEN_706; // @[Multiplier.scala 64:55]
  assign _GEN_708 = 11'h2c4 == fractionSum[12:2] ? 10'h19d : _GEN_707; // @[Multiplier.scala 64:55]
  assign _GEN_709 = 11'h2c5 == fractionSum[12:2] ? 10'h19e : _GEN_708; // @[Multiplier.scala 64:55]
  assign _GEN_710 = 11'h2c6 == fractionSum[12:2] ? 10'h19e : _GEN_709; // @[Multiplier.scala 64:55]
  assign _GEN_711 = 11'h2c7 == fractionSum[12:2] ? 10'h19e : _GEN_710; // @[Multiplier.scala 64:55]
  assign _GEN_712 = 11'h2c8 == fractionSum[12:2] ? 10'h19f : _GEN_711; // @[Multiplier.scala 64:55]
  assign _GEN_713 = 11'h2c9 == fractionSum[12:2] ? 10'h19f : _GEN_712; // @[Multiplier.scala 64:55]
  assign _GEN_714 = 11'h2ca == fractionSum[12:2] ? 10'h19f : _GEN_713; // @[Multiplier.scala 64:55]
  assign _GEN_715 = 11'h2cb == fractionSum[12:2] ? 10'h19f : _GEN_714; // @[Multiplier.scala 64:55]
  assign _GEN_716 = 11'h2cc == fractionSum[12:2] ? 10'h1a0 : _GEN_715; // @[Multiplier.scala 64:55]
  assign _GEN_717 = 11'h2cd == fractionSum[12:2] ? 10'h1a0 : _GEN_716; // @[Multiplier.scala 64:55]
  assign _GEN_718 = 11'h2ce == fractionSum[12:2] ? 10'h1a0 : _GEN_717; // @[Multiplier.scala 64:55]
  assign _GEN_719 = 11'h2cf == fractionSum[12:2] ? 10'h1a0 : _GEN_718; // @[Multiplier.scala 64:55]
  assign _GEN_720 = 11'h2d0 == fractionSum[12:2] ? 10'h1a1 : _GEN_719; // @[Multiplier.scala 64:55]
  assign _GEN_721 = 11'h2d1 == fractionSum[12:2] ? 10'h1a1 : _GEN_720; // @[Multiplier.scala 64:55]
  assign _GEN_722 = 11'h2d2 == fractionSum[12:2] ? 10'h1a1 : _GEN_721; // @[Multiplier.scala 64:55]
  assign _GEN_723 = 11'h2d3 == fractionSum[12:2] ? 10'h1a2 : _GEN_722; // @[Multiplier.scala 64:55]
  assign _GEN_724 = 11'h2d4 == fractionSum[12:2] ? 10'h1a2 : _GEN_723; // @[Multiplier.scala 64:55]
  assign _GEN_725 = 11'h2d5 == fractionSum[12:2] ? 10'h1a2 : _GEN_724; // @[Multiplier.scala 64:55]
  assign _GEN_726 = 11'h2d6 == fractionSum[12:2] ? 10'h1a2 : _GEN_725; // @[Multiplier.scala 64:55]
  assign _GEN_727 = 11'h2d7 == fractionSum[12:2] ? 10'h1a3 : _GEN_726; // @[Multiplier.scala 64:55]
  assign _GEN_728 = 11'h2d8 == fractionSum[12:2] ? 10'h1a3 : _GEN_727; // @[Multiplier.scala 64:55]
  assign _GEN_729 = 11'h2d9 == fractionSum[12:2] ? 10'h1a3 : _GEN_728; // @[Multiplier.scala 64:55]
  assign _GEN_730 = 11'h2da == fractionSum[12:2] ? 10'h1a4 : _GEN_729; // @[Multiplier.scala 64:55]
  assign _GEN_731 = 11'h2db == fractionSum[12:2] ? 10'h1a4 : _GEN_730; // @[Multiplier.scala 64:55]
  assign _GEN_732 = 11'h2dc == fractionSum[12:2] ? 10'h1a4 : _GEN_731; // @[Multiplier.scala 64:55]
  assign _GEN_733 = 11'h2dd == fractionSum[12:2] ? 10'h1a4 : _GEN_732; // @[Multiplier.scala 64:55]
  assign _GEN_734 = 11'h2de == fractionSum[12:2] ? 10'h1a5 : _GEN_733; // @[Multiplier.scala 64:55]
  assign _GEN_735 = 11'h2df == fractionSum[12:2] ? 10'h1a5 : _GEN_734; // @[Multiplier.scala 64:55]
  assign _GEN_736 = 11'h2e0 == fractionSum[12:2] ? 10'h1a5 : _GEN_735; // @[Multiplier.scala 64:55]
  assign _GEN_737 = 11'h2e1 == fractionSum[12:2] ? 10'h1a6 : _GEN_736; // @[Multiplier.scala 64:55]
  assign _GEN_738 = 11'h2e2 == fractionSum[12:2] ? 10'h1a6 : _GEN_737; // @[Multiplier.scala 64:55]
  assign _GEN_739 = 11'h2e3 == fractionSum[12:2] ? 10'h1a6 : _GEN_738; // @[Multiplier.scala 64:55]
  assign _GEN_740 = 11'h2e4 == fractionSum[12:2] ? 10'h1a6 : _GEN_739; // @[Multiplier.scala 64:55]
  assign _GEN_741 = 11'h2e5 == fractionSum[12:2] ? 10'h1a7 : _GEN_740; // @[Multiplier.scala 64:55]
  assign _GEN_742 = 11'h2e6 == fractionSum[12:2] ? 10'h1a7 : _GEN_741; // @[Multiplier.scala 64:55]
  assign _GEN_743 = 11'h2e7 == fractionSum[12:2] ? 10'h1a7 : _GEN_742; // @[Multiplier.scala 64:55]
  assign _GEN_744 = 11'h2e8 == fractionSum[12:2] ? 10'h1a8 : _GEN_743; // @[Multiplier.scala 64:55]
  assign _GEN_745 = 11'h2e9 == fractionSum[12:2] ? 10'h1a8 : _GEN_744; // @[Multiplier.scala 64:55]
  assign _GEN_746 = 11'h2ea == fractionSum[12:2] ? 10'h1a8 : _GEN_745; // @[Multiplier.scala 64:55]
  assign _GEN_747 = 11'h2eb == fractionSum[12:2] ? 10'h1a8 : _GEN_746; // @[Multiplier.scala 64:55]
  assign _GEN_748 = 11'h2ec == fractionSum[12:2] ? 10'h1a9 : _GEN_747; // @[Multiplier.scala 64:55]
  assign _GEN_749 = 11'h2ed == fractionSum[12:2] ? 10'h1a9 : _GEN_748; // @[Multiplier.scala 64:55]
  assign _GEN_750 = 11'h2ee == fractionSum[12:2] ? 10'h1a9 : _GEN_749; // @[Multiplier.scala 64:55]
  assign _GEN_751 = 11'h2ef == fractionSum[12:2] ? 10'h1aa : _GEN_750; // @[Multiplier.scala 64:55]
  assign _GEN_752 = 11'h2f0 == fractionSum[12:2] ? 10'h1aa : _GEN_751; // @[Multiplier.scala 64:55]
  assign _GEN_753 = 11'h2f1 == fractionSum[12:2] ? 10'h1aa : _GEN_752; // @[Multiplier.scala 64:55]
  assign _GEN_754 = 11'h2f2 == fractionSum[12:2] ? 10'h1aa : _GEN_753; // @[Multiplier.scala 64:55]
  assign _GEN_755 = 11'h2f3 == fractionSum[12:2] ? 10'h1ab : _GEN_754; // @[Multiplier.scala 64:55]
  assign _GEN_756 = 11'h2f4 == fractionSum[12:2] ? 10'h1ab : _GEN_755; // @[Multiplier.scala 64:55]
  assign _GEN_757 = 11'h2f5 == fractionSum[12:2] ? 10'h1ab : _GEN_756; // @[Multiplier.scala 64:55]
  assign _GEN_758 = 11'h2f6 == fractionSum[12:2] ? 10'h1ac : _GEN_757; // @[Multiplier.scala 64:55]
  assign _GEN_759 = 11'h2f7 == fractionSum[12:2] ? 10'h1ac : _GEN_758; // @[Multiplier.scala 64:55]
  assign _GEN_760 = 11'h2f8 == fractionSum[12:2] ? 10'h1ac : _GEN_759; // @[Multiplier.scala 64:55]
  assign _GEN_761 = 11'h2f9 == fractionSum[12:2] ? 10'h1ad : _GEN_760; // @[Multiplier.scala 64:55]
  assign _GEN_762 = 11'h2fa == fractionSum[12:2] ? 10'h1ad : _GEN_761; // @[Multiplier.scala 64:55]
  assign _GEN_763 = 11'h2fb == fractionSum[12:2] ? 10'h1ad : _GEN_762; // @[Multiplier.scala 64:55]
  assign _GEN_764 = 11'h2fc == fractionSum[12:2] ? 10'h1ad : _GEN_763; // @[Multiplier.scala 64:55]
  assign _GEN_765 = 11'h2fd == fractionSum[12:2] ? 10'h1ae : _GEN_764; // @[Multiplier.scala 64:55]
  assign _GEN_766 = 11'h2fe == fractionSum[12:2] ? 10'h1ae : _GEN_765; // @[Multiplier.scala 64:55]
  assign _GEN_767 = 11'h2ff == fractionSum[12:2] ? 10'h1ae : _GEN_766; // @[Multiplier.scala 64:55]
  assign _GEN_768 = 11'h300 == fractionSum[12:2] ? 10'h1af : _GEN_767; // @[Multiplier.scala 64:55]
  assign _GEN_769 = 11'h301 == fractionSum[12:2] ? 10'h1af : _GEN_768; // @[Multiplier.scala 64:55]
  assign _GEN_770 = 11'h302 == fractionSum[12:2] ? 10'h1af : _GEN_769; // @[Multiplier.scala 64:55]
  assign _GEN_771 = 11'h303 == fractionSum[12:2] ? 10'h1af : _GEN_770; // @[Multiplier.scala 64:55]
  assign _GEN_772 = 11'h304 == fractionSum[12:2] ? 10'h1b0 : _GEN_771; // @[Multiplier.scala 64:55]
  assign _GEN_773 = 11'h305 == fractionSum[12:2] ? 10'h1b0 : _GEN_772; // @[Multiplier.scala 64:55]
  assign _GEN_774 = 11'h306 == fractionSum[12:2] ? 10'h1b0 : _GEN_773; // @[Multiplier.scala 64:55]
  assign _GEN_775 = 11'h307 == fractionSum[12:2] ? 10'h1b1 : _GEN_774; // @[Multiplier.scala 64:55]
  assign _GEN_776 = 11'h308 == fractionSum[12:2] ? 10'h1b1 : _GEN_775; // @[Multiplier.scala 64:55]
  assign _GEN_777 = 11'h309 == fractionSum[12:2] ? 10'h1b1 : _GEN_776; // @[Multiplier.scala 64:55]
  assign _GEN_778 = 11'h30a == fractionSum[12:2] ? 10'h1b1 : _GEN_777; // @[Multiplier.scala 64:55]
  assign _GEN_779 = 11'h30b == fractionSum[12:2] ? 10'h1b2 : _GEN_778; // @[Multiplier.scala 64:55]
  assign _GEN_780 = 11'h30c == fractionSum[12:2] ? 10'h1b2 : _GEN_779; // @[Multiplier.scala 64:55]
  assign _GEN_781 = 11'h30d == fractionSum[12:2] ? 10'h1b2 : _GEN_780; // @[Multiplier.scala 64:55]
  assign _GEN_782 = 11'h30e == fractionSum[12:2] ? 10'h1b3 : _GEN_781; // @[Multiplier.scala 64:55]
  assign _GEN_783 = 11'h30f == fractionSum[12:2] ? 10'h1b3 : _GEN_782; // @[Multiplier.scala 64:55]
  assign _GEN_784 = 11'h310 == fractionSum[12:2] ? 10'h1b3 : _GEN_783; // @[Multiplier.scala 64:55]
  assign _GEN_785 = 11'h311 == fractionSum[12:2] ? 10'h1b4 : _GEN_784; // @[Multiplier.scala 64:55]
  assign _GEN_786 = 11'h312 == fractionSum[12:2] ? 10'h1b4 : _GEN_785; // @[Multiplier.scala 64:55]
  assign _GEN_787 = 11'h313 == fractionSum[12:2] ? 10'h1b4 : _GEN_786; // @[Multiplier.scala 64:55]
  assign _GEN_788 = 11'h314 == fractionSum[12:2] ? 10'h1b4 : _GEN_787; // @[Multiplier.scala 64:55]
  assign _GEN_789 = 11'h315 == fractionSum[12:2] ? 10'h1b5 : _GEN_788; // @[Multiplier.scala 64:55]
  assign _GEN_790 = 11'h316 == fractionSum[12:2] ? 10'h1b5 : _GEN_789; // @[Multiplier.scala 64:55]
  assign _GEN_791 = 11'h317 == fractionSum[12:2] ? 10'h1b5 : _GEN_790; // @[Multiplier.scala 64:55]
  assign _GEN_792 = 11'h318 == fractionSum[12:2] ? 10'h1b6 : _GEN_791; // @[Multiplier.scala 64:55]
  assign _GEN_793 = 11'h319 == fractionSum[12:2] ? 10'h1b6 : _GEN_792; // @[Multiplier.scala 64:55]
  assign _GEN_794 = 11'h31a == fractionSum[12:2] ? 10'h1b6 : _GEN_793; // @[Multiplier.scala 64:55]
  assign _GEN_795 = 11'h31b == fractionSum[12:2] ? 10'h1b6 : _GEN_794; // @[Multiplier.scala 64:55]
  assign _GEN_796 = 11'h31c == fractionSum[12:2] ? 10'h1b7 : _GEN_795; // @[Multiplier.scala 64:55]
  assign _GEN_797 = 11'h31d == fractionSum[12:2] ? 10'h1b7 : _GEN_796; // @[Multiplier.scala 64:55]
  assign _GEN_798 = 11'h31e == fractionSum[12:2] ? 10'h1b7 : _GEN_797; // @[Multiplier.scala 64:55]
  assign _GEN_799 = 11'h31f == fractionSum[12:2] ? 10'h1b8 : _GEN_798; // @[Multiplier.scala 64:55]
  assign _GEN_800 = 11'h320 == fractionSum[12:2] ? 10'h1b8 : _GEN_799; // @[Multiplier.scala 64:55]
  assign _GEN_801 = 11'h321 == fractionSum[12:2] ? 10'h1b8 : _GEN_800; // @[Multiplier.scala 64:55]
  assign _GEN_802 = 11'h322 == fractionSum[12:2] ? 10'h1b9 : _GEN_801; // @[Multiplier.scala 64:55]
  assign _GEN_803 = 11'h323 == fractionSum[12:2] ? 10'h1b9 : _GEN_802; // @[Multiplier.scala 64:55]
  assign _GEN_804 = 11'h324 == fractionSum[12:2] ? 10'h1b9 : _GEN_803; // @[Multiplier.scala 64:55]
  assign _GEN_805 = 11'h325 == fractionSum[12:2] ? 10'h1b9 : _GEN_804; // @[Multiplier.scala 64:55]
  assign _GEN_806 = 11'h326 == fractionSum[12:2] ? 10'h1ba : _GEN_805; // @[Multiplier.scala 64:55]
  assign _GEN_807 = 11'h327 == fractionSum[12:2] ? 10'h1ba : _GEN_806; // @[Multiplier.scala 64:55]
  assign _GEN_808 = 11'h328 == fractionSum[12:2] ? 10'h1ba : _GEN_807; // @[Multiplier.scala 64:55]
  assign _GEN_809 = 11'h329 == fractionSum[12:2] ? 10'h1bb : _GEN_808; // @[Multiplier.scala 64:55]
  assign _GEN_810 = 11'h32a == fractionSum[12:2] ? 10'h1bb : _GEN_809; // @[Multiplier.scala 64:55]
  assign _GEN_811 = 11'h32b == fractionSum[12:2] ? 10'h1bb : _GEN_810; // @[Multiplier.scala 64:55]
  assign _GEN_812 = 11'h32c == fractionSum[12:2] ? 10'h1bc : _GEN_811; // @[Multiplier.scala 64:55]
  assign _GEN_813 = 11'h32d == fractionSum[12:2] ? 10'h1bc : _GEN_812; // @[Multiplier.scala 64:55]
  assign _GEN_814 = 11'h32e == fractionSum[12:2] ? 10'h1bc : _GEN_813; // @[Multiplier.scala 64:55]
  assign _GEN_815 = 11'h32f == fractionSum[12:2] ? 10'h1bc : _GEN_814; // @[Multiplier.scala 64:55]
  assign _GEN_816 = 11'h330 == fractionSum[12:2] ? 10'h1bd : _GEN_815; // @[Multiplier.scala 64:55]
  assign _GEN_817 = 11'h331 == fractionSum[12:2] ? 10'h1bd : _GEN_816; // @[Multiplier.scala 64:55]
  assign _GEN_818 = 11'h332 == fractionSum[12:2] ? 10'h1bd : _GEN_817; // @[Multiplier.scala 64:55]
  assign _GEN_819 = 11'h333 == fractionSum[12:2] ? 10'h1be : _GEN_818; // @[Multiplier.scala 64:55]
  assign _GEN_820 = 11'h334 == fractionSum[12:2] ? 10'h1be : _GEN_819; // @[Multiplier.scala 64:55]
  assign _GEN_821 = 11'h335 == fractionSum[12:2] ? 10'h1be : _GEN_820; // @[Multiplier.scala 64:55]
  assign _GEN_822 = 11'h336 == fractionSum[12:2] ? 10'h1bf : _GEN_821; // @[Multiplier.scala 64:55]
  assign _GEN_823 = 11'h337 == fractionSum[12:2] ? 10'h1bf : _GEN_822; // @[Multiplier.scala 64:55]
  assign _GEN_824 = 11'h338 == fractionSum[12:2] ? 10'h1bf : _GEN_823; // @[Multiplier.scala 64:55]
  assign _GEN_825 = 11'h339 == fractionSum[12:2] ? 10'h1bf : _GEN_824; // @[Multiplier.scala 64:55]
  assign _GEN_826 = 11'h33a == fractionSum[12:2] ? 10'h1c0 : _GEN_825; // @[Multiplier.scala 64:55]
  assign _GEN_827 = 11'h33b == fractionSum[12:2] ? 10'h1c0 : _GEN_826; // @[Multiplier.scala 64:55]
  assign _GEN_828 = 11'h33c == fractionSum[12:2] ? 10'h1c0 : _GEN_827; // @[Multiplier.scala 64:55]
  assign _GEN_829 = 11'h33d == fractionSum[12:2] ? 10'h1c1 : _GEN_828; // @[Multiplier.scala 64:55]
  assign _GEN_830 = 11'h33e == fractionSum[12:2] ? 10'h1c1 : _GEN_829; // @[Multiplier.scala 64:55]
  assign _GEN_831 = 11'h33f == fractionSum[12:2] ? 10'h1c1 : _GEN_830; // @[Multiplier.scala 64:55]
  assign _GEN_832 = 11'h340 == fractionSum[12:2] ? 10'h1c2 : _GEN_831; // @[Multiplier.scala 64:55]
  assign _GEN_833 = 11'h341 == fractionSum[12:2] ? 10'h1c2 : _GEN_832; // @[Multiplier.scala 64:55]
  assign _GEN_834 = 11'h342 == fractionSum[12:2] ? 10'h1c2 : _GEN_833; // @[Multiplier.scala 64:55]
  assign _GEN_835 = 11'h343 == fractionSum[12:2] ? 10'h1c3 : _GEN_834; // @[Multiplier.scala 64:55]
  assign _GEN_836 = 11'h344 == fractionSum[12:2] ? 10'h1c3 : _GEN_835; // @[Multiplier.scala 64:55]
  assign _GEN_837 = 11'h345 == fractionSum[12:2] ? 10'h1c3 : _GEN_836; // @[Multiplier.scala 64:55]
  assign _GEN_838 = 11'h346 == fractionSum[12:2] ? 10'h1c3 : _GEN_837; // @[Multiplier.scala 64:55]
  assign _GEN_839 = 11'h347 == fractionSum[12:2] ? 10'h1c4 : _GEN_838; // @[Multiplier.scala 64:55]
  assign _GEN_840 = 11'h348 == fractionSum[12:2] ? 10'h1c4 : _GEN_839; // @[Multiplier.scala 64:55]
  assign _GEN_841 = 11'h349 == fractionSum[12:2] ? 10'h1c4 : _GEN_840; // @[Multiplier.scala 64:55]
  assign _GEN_842 = 11'h34a == fractionSum[12:2] ? 10'h1c5 : _GEN_841; // @[Multiplier.scala 64:55]
  assign _GEN_843 = 11'h34b == fractionSum[12:2] ? 10'h1c5 : _GEN_842; // @[Multiplier.scala 64:55]
  assign _GEN_844 = 11'h34c == fractionSum[12:2] ? 10'h1c5 : _GEN_843; // @[Multiplier.scala 64:55]
  assign _GEN_845 = 11'h34d == fractionSum[12:2] ? 10'h1c6 : _GEN_844; // @[Multiplier.scala 64:55]
  assign _GEN_846 = 11'h34e == fractionSum[12:2] ? 10'h1c6 : _GEN_845; // @[Multiplier.scala 64:55]
  assign _GEN_847 = 11'h34f == fractionSum[12:2] ? 10'h1c6 : _GEN_846; // @[Multiplier.scala 64:55]
  assign _GEN_848 = 11'h350 == fractionSum[12:2] ? 10'h1c6 : _GEN_847; // @[Multiplier.scala 64:55]
  assign _GEN_849 = 11'h351 == fractionSum[12:2] ? 10'h1c7 : _GEN_848; // @[Multiplier.scala 64:55]
  assign _GEN_850 = 11'h352 == fractionSum[12:2] ? 10'h1c7 : _GEN_849; // @[Multiplier.scala 64:55]
  assign _GEN_851 = 11'h353 == fractionSum[12:2] ? 10'h1c7 : _GEN_850; // @[Multiplier.scala 64:55]
  assign _GEN_852 = 11'h354 == fractionSum[12:2] ? 10'h1c8 : _GEN_851; // @[Multiplier.scala 64:55]
  assign _GEN_853 = 11'h355 == fractionSum[12:2] ? 10'h1c8 : _GEN_852; // @[Multiplier.scala 64:55]
  assign _GEN_854 = 11'h356 == fractionSum[12:2] ? 10'h1c8 : _GEN_853; // @[Multiplier.scala 64:55]
  assign _GEN_855 = 11'h357 == fractionSum[12:2] ? 10'h1c9 : _GEN_854; // @[Multiplier.scala 64:55]
  assign _GEN_856 = 11'h358 == fractionSum[12:2] ? 10'h1c9 : _GEN_855; // @[Multiplier.scala 64:55]
  assign _GEN_857 = 11'h359 == fractionSum[12:2] ? 10'h1c9 : _GEN_856; // @[Multiplier.scala 64:55]
  assign _GEN_858 = 11'h35a == fractionSum[12:2] ? 10'h1ca : _GEN_857; // @[Multiplier.scala 64:55]
  assign _GEN_859 = 11'h35b == fractionSum[12:2] ? 10'h1ca : _GEN_858; // @[Multiplier.scala 64:55]
  assign _GEN_860 = 11'h35c == fractionSum[12:2] ? 10'h1ca : _GEN_859; // @[Multiplier.scala 64:55]
  assign _GEN_861 = 11'h35d == fractionSum[12:2] ? 10'h1cb : _GEN_860; // @[Multiplier.scala 64:55]
  assign _GEN_862 = 11'h35e == fractionSum[12:2] ? 10'h1cb : _GEN_861; // @[Multiplier.scala 64:55]
  assign _GEN_863 = 11'h35f == fractionSum[12:2] ? 10'h1cb : _GEN_862; // @[Multiplier.scala 64:55]
  assign _GEN_864 = 11'h360 == fractionSum[12:2] ? 10'h1cb : _GEN_863; // @[Multiplier.scala 64:55]
  assign _GEN_865 = 11'h361 == fractionSum[12:2] ? 10'h1cc : _GEN_864; // @[Multiplier.scala 64:55]
  assign _GEN_866 = 11'h362 == fractionSum[12:2] ? 10'h1cc : _GEN_865; // @[Multiplier.scala 64:55]
  assign _GEN_867 = 11'h363 == fractionSum[12:2] ? 10'h1cc : _GEN_866; // @[Multiplier.scala 64:55]
  assign _GEN_868 = 11'h364 == fractionSum[12:2] ? 10'h1cd : _GEN_867; // @[Multiplier.scala 64:55]
  assign _GEN_869 = 11'h365 == fractionSum[12:2] ? 10'h1cd : _GEN_868; // @[Multiplier.scala 64:55]
  assign _GEN_870 = 11'h366 == fractionSum[12:2] ? 10'h1cd : _GEN_869; // @[Multiplier.scala 64:55]
  assign _GEN_871 = 11'h367 == fractionSum[12:2] ? 10'h1ce : _GEN_870; // @[Multiplier.scala 64:55]
  assign _GEN_872 = 11'h368 == fractionSum[12:2] ? 10'h1ce : _GEN_871; // @[Multiplier.scala 64:55]
  assign _GEN_873 = 11'h369 == fractionSum[12:2] ? 10'h1ce : _GEN_872; // @[Multiplier.scala 64:55]
  assign _GEN_874 = 11'h36a == fractionSum[12:2] ? 10'h1cf : _GEN_873; // @[Multiplier.scala 64:55]
  assign _GEN_875 = 11'h36b == fractionSum[12:2] ? 10'h1cf : _GEN_874; // @[Multiplier.scala 64:55]
  assign _GEN_876 = 11'h36c == fractionSum[12:2] ? 10'h1cf : _GEN_875; // @[Multiplier.scala 64:55]
  assign _GEN_877 = 11'h36d == fractionSum[12:2] ? 10'h1d0 : _GEN_876; // @[Multiplier.scala 64:55]
  assign _GEN_878 = 11'h36e == fractionSum[12:2] ? 10'h1d0 : _GEN_877; // @[Multiplier.scala 64:55]
  assign _GEN_879 = 11'h36f == fractionSum[12:2] ? 10'h1d0 : _GEN_878; // @[Multiplier.scala 64:55]
  assign _GEN_880 = 11'h370 == fractionSum[12:2] ? 10'h1d0 : _GEN_879; // @[Multiplier.scala 64:55]
  assign _GEN_881 = 11'h371 == fractionSum[12:2] ? 10'h1d1 : _GEN_880; // @[Multiplier.scala 64:55]
  assign _GEN_882 = 11'h372 == fractionSum[12:2] ? 10'h1d1 : _GEN_881; // @[Multiplier.scala 64:55]
  assign _GEN_883 = 11'h373 == fractionSum[12:2] ? 10'h1d1 : _GEN_882; // @[Multiplier.scala 64:55]
  assign _GEN_884 = 11'h374 == fractionSum[12:2] ? 10'h1d2 : _GEN_883; // @[Multiplier.scala 64:55]
  assign _GEN_885 = 11'h375 == fractionSum[12:2] ? 10'h1d2 : _GEN_884; // @[Multiplier.scala 64:55]
  assign _GEN_886 = 11'h376 == fractionSum[12:2] ? 10'h1d2 : _GEN_885; // @[Multiplier.scala 64:55]
  assign _GEN_887 = 11'h377 == fractionSum[12:2] ? 10'h1d3 : _GEN_886; // @[Multiplier.scala 64:55]
  assign _GEN_888 = 11'h378 == fractionSum[12:2] ? 10'h1d3 : _GEN_887; // @[Multiplier.scala 64:55]
  assign _GEN_889 = 11'h379 == fractionSum[12:2] ? 10'h1d3 : _GEN_888; // @[Multiplier.scala 64:55]
  assign _GEN_890 = 11'h37a == fractionSum[12:2] ? 10'h1d4 : _GEN_889; // @[Multiplier.scala 64:55]
  assign _GEN_891 = 11'h37b == fractionSum[12:2] ? 10'h1d4 : _GEN_890; // @[Multiplier.scala 64:55]
  assign _GEN_892 = 11'h37c == fractionSum[12:2] ? 10'h1d4 : _GEN_891; // @[Multiplier.scala 64:55]
  assign _GEN_893 = 11'h37d == fractionSum[12:2] ? 10'h1d5 : _GEN_892; // @[Multiplier.scala 64:55]
  assign _GEN_894 = 11'h37e == fractionSum[12:2] ? 10'h1d5 : _GEN_893; // @[Multiplier.scala 64:55]
  assign _GEN_895 = 11'h37f == fractionSum[12:2] ? 10'h1d5 : _GEN_894; // @[Multiplier.scala 64:55]
  assign _GEN_896 = 11'h380 == fractionSum[12:2] ? 10'h1d6 : _GEN_895; // @[Multiplier.scala 64:55]
  assign _GEN_897 = 11'h381 == fractionSum[12:2] ? 10'h1d6 : _GEN_896; // @[Multiplier.scala 64:55]
  assign _GEN_898 = 11'h382 == fractionSum[12:2] ? 10'h1d6 : _GEN_897; // @[Multiplier.scala 64:55]
  assign _GEN_899 = 11'h383 == fractionSum[12:2] ? 10'h1d6 : _GEN_898; // @[Multiplier.scala 64:55]
  assign _GEN_900 = 11'h384 == fractionSum[12:2] ? 10'h1d7 : _GEN_899; // @[Multiplier.scala 64:55]
  assign _GEN_901 = 11'h385 == fractionSum[12:2] ? 10'h1d7 : _GEN_900; // @[Multiplier.scala 64:55]
  assign _GEN_902 = 11'h386 == fractionSum[12:2] ? 10'h1d7 : _GEN_901; // @[Multiplier.scala 64:55]
  assign _GEN_903 = 11'h387 == fractionSum[12:2] ? 10'h1d8 : _GEN_902; // @[Multiplier.scala 64:55]
  assign _GEN_904 = 11'h388 == fractionSum[12:2] ? 10'h1d8 : _GEN_903; // @[Multiplier.scala 64:55]
  assign _GEN_905 = 11'h389 == fractionSum[12:2] ? 10'h1d8 : _GEN_904; // @[Multiplier.scala 64:55]
  assign _GEN_906 = 11'h38a == fractionSum[12:2] ? 10'h1d9 : _GEN_905; // @[Multiplier.scala 64:55]
  assign _GEN_907 = 11'h38b == fractionSum[12:2] ? 10'h1d9 : _GEN_906; // @[Multiplier.scala 64:55]
  assign _GEN_908 = 11'h38c == fractionSum[12:2] ? 10'h1d9 : _GEN_907; // @[Multiplier.scala 64:55]
  assign _GEN_909 = 11'h38d == fractionSum[12:2] ? 10'h1da : _GEN_908; // @[Multiplier.scala 64:55]
  assign _GEN_910 = 11'h38e == fractionSum[12:2] ? 10'h1da : _GEN_909; // @[Multiplier.scala 64:55]
  assign _GEN_911 = 11'h38f == fractionSum[12:2] ? 10'h1da : _GEN_910; // @[Multiplier.scala 64:55]
  assign _GEN_912 = 11'h390 == fractionSum[12:2] ? 10'h1db : _GEN_911; // @[Multiplier.scala 64:55]
  assign _GEN_913 = 11'h391 == fractionSum[12:2] ? 10'h1db : _GEN_912; // @[Multiplier.scala 64:55]
  assign _GEN_914 = 11'h392 == fractionSum[12:2] ? 10'h1db : _GEN_913; // @[Multiplier.scala 64:55]
  assign _GEN_915 = 11'h393 == fractionSum[12:2] ? 10'h1dc : _GEN_914; // @[Multiplier.scala 64:55]
  assign _GEN_916 = 11'h394 == fractionSum[12:2] ? 10'h1dc : _GEN_915; // @[Multiplier.scala 64:55]
  assign _GEN_917 = 11'h395 == fractionSum[12:2] ? 10'h1dc : _GEN_916; // @[Multiplier.scala 64:55]
  assign _GEN_918 = 11'h396 == fractionSum[12:2] ? 10'h1dd : _GEN_917; // @[Multiplier.scala 64:55]
  assign _GEN_919 = 11'h397 == fractionSum[12:2] ? 10'h1dd : _GEN_918; // @[Multiplier.scala 64:55]
  assign _GEN_920 = 11'h398 == fractionSum[12:2] ? 10'h1dd : _GEN_919; // @[Multiplier.scala 64:55]
  assign _GEN_921 = 11'h399 == fractionSum[12:2] ? 10'h1de : _GEN_920; // @[Multiplier.scala 64:55]
  assign _GEN_922 = 11'h39a == fractionSum[12:2] ? 10'h1de : _GEN_921; // @[Multiplier.scala 64:55]
  assign _GEN_923 = 11'h39b == fractionSum[12:2] ? 10'h1de : _GEN_922; // @[Multiplier.scala 64:55]
  assign _GEN_924 = 11'h39c == fractionSum[12:2] ? 10'h1de : _GEN_923; // @[Multiplier.scala 64:55]
  assign _GEN_925 = 11'h39d == fractionSum[12:2] ? 10'h1df : _GEN_924; // @[Multiplier.scala 64:55]
  assign _GEN_926 = 11'h39e == fractionSum[12:2] ? 10'h1df : _GEN_925; // @[Multiplier.scala 64:55]
  assign _GEN_927 = 11'h39f == fractionSum[12:2] ? 10'h1df : _GEN_926; // @[Multiplier.scala 64:55]
  assign _GEN_928 = 11'h3a0 == fractionSum[12:2] ? 10'h1e0 : _GEN_927; // @[Multiplier.scala 64:55]
  assign _GEN_929 = 11'h3a1 == fractionSum[12:2] ? 10'h1e0 : _GEN_928; // @[Multiplier.scala 64:55]
  assign _GEN_930 = 11'h3a2 == fractionSum[12:2] ? 10'h1e0 : _GEN_929; // @[Multiplier.scala 64:55]
  assign _GEN_931 = 11'h3a3 == fractionSum[12:2] ? 10'h1e1 : _GEN_930; // @[Multiplier.scala 64:55]
  assign _GEN_932 = 11'h3a4 == fractionSum[12:2] ? 10'h1e1 : _GEN_931; // @[Multiplier.scala 64:55]
  assign _GEN_933 = 11'h3a5 == fractionSum[12:2] ? 10'h1e1 : _GEN_932; // @[Multiplier.scala 64:55]
  assign _GEN_934 = 11'h3a6 == fractionSum[12:2] ? 10'h1e2 : _GEN_933; // @[Multiplier.scala 64:55]
  assign _GEN_935 = 11'h3a7 == fractionSum[12:2] ? 10'h1e2 : _GEN_934; // @[Multiplier.scala 64:55]
  assign _GEN_936 = 11'h3a8 == fractionSum[12:2] ? 10'h1e2 : _GEN_935; // @[Multiplier.scala 64:55]
  assign _GEN_937 = 11'h3a9 == fractionSum[12:2] ? 10'h1e3 : _GEN_936; // @[Multiplier.scala 64:55]
  assign _GEN_938 = 11'h3aa == fractionSum[12:2] ? 10'h1e3 : _GEN_937; // @[Multiplier.scala 64:55]
  assign _GEN_939 = 11'h3ab == fractionSum[12:2] ? 10'h1e3 : _GEN_938; // @[Multiplier.scala 64:55]
  assign _GEN_940 = 11'h3ac == fractionSum[12:2] ? 10'h1e4 : _GEN_939; // @[Multiplier.scala 64:55]
  assign _GEN_941 = 11'h3ad == fractionSum[12:2] ? 10'h1e4 : _GEN_940; // @[Multiplier.scala 64:55]
  assign _GEN_942 = 11'h3ae == fractionSum[12:2] ? 10'h1e4 : _GEN_941; // @[Multiplier.scala 64:55]
  assign _GEN_943 = 11'h3af == fractionSum[12:2] ? 10'h1e5 : _GEN_942; // @[Multiplier.scala 64:55]
  assign _GEN_944 = 11'h3b0 == fractionSum[12:2] ? 10'h1e5 : _GEN_943; // @[Multiplier.scala 64:55]
  assign _GEN_945 = 11'h3b1 == fractionSum[12:2] ? 10'h1e5 : _GEN_944; // @[Multiplier.scala 64:55]
  assign _GEN_946 = 11'h3b2 == fractionSum[12:2] ? 10'h1e6 : _GEN_945; // @[Multiplier.scala 64:55]
  assign _GEN_947 = 11'h3b3 == fractionSum[12:2] ? 10'h1e6 : _GEN_946; // @[Multiplier.scala 64:55]
  assign _GEN_948 = 11'h3b4 == fractionSum[12:2] ? 10'h1e6 : _GEN_947; // @[Multiplier.scala 64:55]
  assign _GEN_949 = 11'h3b5 == fractionSum[12:2] ? 10'h1e7 : _GEN_948; // @[Multiplier.scala 64:55]
  assign _GEN_950 = 11'h3b6 == fractionSum[12:2] ? 10'h1e7 : _GEN_949; // @[Multiplier.scala 64:55]
  assign _GEN_951 = 11'h3b7 == fractionSum[12:2] ? 10'h1e7 : _GEN_950; // @[Multiplier.scala 64:55]
  assign _GEN_952 = 11'h3b8 == fractionSum[12:2] ? 10'h1e8 : _GEN_951; // @[Multiplier.scala 64:55]
  assign _GEN_953 = 11'h3b9 == fractionSum[12:2] ? 10'h1e8 : _GEN_952; // @[Multiplier.scala 64:55]
  assign _GEN_954 = 11'h3ba == fractionSum[12:2] ? 10'h1e8 : _GEN_953; // @[Multiplier.scala 64:55]
  assign _GEN_955 = 11'h3bb == fractionSum[12:2] ? 10'h1e9 : _GEN_954; // @[Multiplier.scala 64:55]
  assign _GEN_956 = 11'h3bc == fractionSum[12:2] ? 10'h1e9 : _GEN_955; // @[Multiplier.scala 64:55]
  assign _GEN_957 = 11'h3bd == fractionSum[12:2] ? 10'h1e9 : _GEN_956; // @[Multiplier.scala 64:55]
  assign _GEN_958 = 11'h3be == fractionSum[12:2] ? 10'h1ea : _GEN_957; // @[Multiplier.scala 64:55]
  assign _GEN_959 = 11'h3bf == fractionSum[12:2] ? 10'h1ea : _GEN_958; // @[Multiplier.scala 64:55]
  assign _GEN_960 = 11'h3c0 == fractionSum[12:2] ? 10'h1ea : _GEN_959; // @[Multiplier.scala 64:55]
  assign _GEN_961 = 11'h3c1 == fractionSum[12:2] ? 10'h1eb : _GEN_960; // @[Multiplier.scala 64:55]
  assign _GEN_962 = 11'h3c2 == fractionSum[12:2] ? 10'h1eb : _GEN_961; // @[Multiplier.scala 64:55]
  assign _GEN_963 = 11'h3c3 == fractionSum[12:2] ? 10'h1eb : _GEN_962; // @[Multiplier.scala 64:55]
  assign _GEN_964 = 11'h3c4 == fractionSum[12:2] ? 10'h1ec : _GEN_963; // @[Multiplier.scala 64:55]
  assign _GEN_965 = 11'h3c5 == fractionSum[12:2] ? 10'h1ec : _GEN_964; // @[Multiplier.scala 64:55]
  assign _GEN_966 = 11'h3c6 == fractionSum[12:2] ? 10'h1ec : _GEN_965; // @[Multiplier.scala 64:55]
  assign _GEN_967 = 11'h3c7 == fractionSum[12:2] ? 10'h1ed : _GEN_966; // @[Multiplier.scala 64:55]
  assign _GEN_968 = 11'h3c8 == fractionSum[12:2] ? 10'h1ed : _GEN_967; // @[Multiplier.scala 64:55]
  assign _GEN_969 = 11'h3c9 == fractionSum[12:2] ? 10'h1ed : _GEN_968; // @[Multiplier.scala 64:55]
  assign _GEN_970 = 11'h3ca == fractionSum[12:2] ? 10'h1ee : _GEN_969; // @[Multiplier.scala 64:55]
  assign _GEN_971 = 11'h3cb == fractionSum[12:2] ? 10'h1ee : _GEN_970; // @[Multiplier.scala 64:55]
  assign _GEN_972 = 11'h3cc == fractionSum[12:2] ? 10'h1ee : _GEN_971; // @[Multiplier.scala 64:55]
  assign _GEN_973 = 11'h3cd == fractionSum[12:2] ? 10'h1ef : _GEN_972; // @[Multiplier.scala 64:55]
  assign _GEN_974 = 11'h3ce == fractionSum[12:2] ? 10'h1ef : _GEN_973; // @[Multiplier.scala 64:55]
  assign _GEN_975 = 11'h3cf == fractionSum[12:2] ? 10'h1ef : _GEN_974; // @[Multiplier.scala 64:55]
  assign _GEN_976 = 11'h3d0 == fractionSum[12:2] ? 10'h1f0 : _GEN_975; // @[Multiplier.scala 64:55]
  assign _GEN_977 = 11'h3d1 == fractionSum[12:2] ? 10'h1f0 : _GEN_976; // @[Multiplier.scala 64:55]
  assign _GEN_978 = 11'h3d2 == fractionSum[12:2] ? 10'h1f0 : _GEN_977; // @[Multiplier.scala 64:55]
  assign _GEN_979 = 11'h3d3 == fractionSum[12:2] ? 10'h1f1 : _GEN_978; // @[Multiplier.scala 64:55]
  assign _GEN_980 = 11'h3d4 == fractionSum[12:2] ? 10'h1f1 : _GEN_979; // @[Multiplier.scala 64:55]
  assign _GEN_981 = 11'h3d5 == fractionSum[12:2] ? 10'h1f1 : _GEN_980; // @[Multiplier.scala 64:55]
  assign _GEN_982 = 11'h3d6 == fractionSum[12:2] ? 10'h1f2 : _GEN_981; // @[Multiplier.scala 64:55]
  assign _GEN_983 = 11'h3d7 == fractionSum[12:2] ? 10'h1f2 : _GEN_982; // @[Multiplier.scala 64:55]
  assign _GEN_984 = 11'h3d8 == fractionSum[12:2] ? 10'h1f2 : _GEN_983; // @[Multiplier.scala 64:55]
  assign _GEN_985 = 11'h3d9 == fractionSum[12:2] ? 10'h1f3 : _GEN_984; // @[Multiplier.scala 64:55]
  assign _GEN_986 = 11'h3da == fractionSum[12:2] ? 10'h1f3 : _GEN_985; // @[Multiplier.scala 64:55]
  assign _GEN_987 = 11'h3db == fractionSum[12:2] ? 10'h1f3 : _GEN_986; // @[Multiplier.scala 64:55]
  assign _GEN_988 = 11'h3dc == fractionSum[12:2] ? 10'h1f4 : _GEN_987; // @[Multiplier.scala 64:55]
  assign _GEN_989 = 11'h3dd == fractionSum[12:2] ? 10'h1f4 : _GEN_988; // @[Multiplier.scala 64:55]
  assign _GEN_990 = 11'h3de == fractionSum[12:2] ? 10'h1f4 : _GEN_989; // @[Multiplier.scala 64:55]
  assign _GEN_991 = 11'h3df == fractionSum[12:2] ? 10'h1f5 : _GEN_990; // @[Multiplier.scala 64:55]
  assign _GEN_992 = 11'h3e0 == fractionSum[12:2] ? 10'h1f5 : _GEN_991; // @[Multiplier.scala 64:55]
  assign _GEN_993 = 11'h3e1 == fractionSum[12:2] ? 10'h1f5 : _GEN_992; // @[Multiplier.scala 64:55]
  assign _GEN_994 = 11'h3e2 == fractionSum[12:2] ? 10'h1f6 : _GEN_993; // @[Multiplier.scala 64:55]
  assign _GEN_995 = 11'h3e3 == fractionSum[12:2] ? 10'h1f6 : _GEN_994; // @[Multiplier.scala 64:55]
  assign _GEN_996 = 11'h3e4 == fractionSum[12:2] ? 10'h1f6 : _GEN_995; // @[Multiplier.scala 64:55]
  assign _GEN_997 = 11'h3e5 == fractionSum[12:2] ? 10'h1f7 : _GEN_996; // @[Multiplier.scala 64:55]
  assign _GEN_998 = 11'h3e6 == fractionSum[12:2] ? 10'h1f7 : _GEN_997; // @[Multiplier.scala 64:55]
  assign _GEN_999 = 11'h3e7 == fractionSum[12:2] ? 10'h1f7 : _GEN_998; // @[Multiplier.scala 64:55]
  assign _GEN_1000 = 11'h3e8 == fractionSum[12:2] ? 10'h1f8 : _GEN_999; // @[Multiplier.scala 64:55]
  assign _GEN_1001 = 11'h3e9 == fractionSum[12:2] ? 10'h1f8 : _GEN_1000; // @[Multiplier.scala 64:55]
  assign _GEN_1002 = 11'h3ea == fractionSum[12:2] ? 10'h1f8 : _GEN_1001; // @[Multiplier.scala 64:55]
  assign _GEN_1003 = 11'h3eb == fractionSum[12:2] ? 10'h1f9 : _GEN_1002; // @[Multiplier.scala 64:55]
  assign _GEN_1004 = 11'h3ec == fractionSum[12:2] ? 10'h1f9 : _GEN_1003; // @[Multiplier.scala 64:55]
  assign _GEN_1005 = 11'h3ed == fractionSum[12:2] ? 10'h1f9 : _GEN_1004; // @[Multiplier.scala 64:55]
  assign _GEN_1006 = 11'h3ee == fractionSum[12:2] ? 10'h1fa : _GEN_1005; // @[Multiplier.scala 64:55]
  assign _GEN_1007 = 11'h3ef == fractionSum[12:2] ? 10'h1fa : _GEN_1006; // @[Multiplier.scala 64:55]
  assign _GEN_1008 = 11'h3f0 == fractionSum[12:2] ? 10'h1fa : _GEN_1007; // @[Multiplier.scala 64:55]
  assign _GEN_1009 = 11'h3f1 == fractionSum[12:2] ? 10'h1fb : _GEN_1008; // @[Multiplier.scala 64:55]
  assign _GEN_1010 = 11'h3f2 == fractionSum[12:2] ? 10'h1fb : _GEN_1009; // @[Multiplier.scala 64:55]
  assign _GEN_1011 = 11'h3f3 == fractionSum[12:2] ? 10'h1fc : _GEN_1010; // @[Multiplier.scala 64:55]
  assign _GEN_1012 = 11'h3f4 == fractionSum[12:2] ? 10'h1fc : _GEN_1011; // @[Multiplier.scala 64:55]
  assign _GEN_1013 = 11'h3f5 == fractionSum[12:2] ? 10'h1fc : _GEN_1012; // @[Multiplier.scala 64:55]
  assign _GEN_1014 = 11'h3f6 == fractionSum[12:2] ? 10'h1fd : _GEN_1013; // @[Multiplier.scala 64:55]
  assign _GEN_1015 = 11'h3f7 == fractionSum[12:2] ? 10'h1fd : _GEN_1014; // @[Multiplier.scala 64:55]
  assign _GEN_1016 = 11'h3f8 == fractionSum[12:2] ? 10'h1fd : _GEN_1015; // @[Multiplier.scala 64:55]
  assign _GEN_1017 = 11'h3f9 == fractionSum[12:2] ? 10'h1fe : _GEN_1016; // @[Multiplier.scala 64:55]
  assign _GEN_1018 = 11'h3fa == fractionSum[12:2] ? 10'h1fe : _GEN_1017; // @[Multiplier.scala 64:55]
  assign _GEN_1019 = 11'h3fb == fractionSum[12:2] ? 10'h1fe : _GEN_1018; // @[Multiplier.scala 64:55]
  assign _GEN_1020 = 11'h3fc == fractionSum[12:2] ? 10'h1ff : _GEN_1019; // @[Multiplier.scala 64:55]
  assign _GEN_1021 = 11'h3fd == fractionSum[12:2] ? 10'h1ff : _GEN_1020; // @[Multiplier.scala 64:55]
  assign _GEN_1022 = 11'h3fe == fractionSum[12:2] ? 10'h1ff : _GEN_1021; // @[Multiplier.scala 64:55]
  assign _GEN_1023 = 11'h3ff == fractionSum[12:2] ? 10'h200 : _GEN_1022; // @[Multiplier.scala 64:55]
  assign _GEN_1024 = 11'h400 == fractionSum[12:2] ? 10'h200 : _GEN_1023; // @[Multiplier.scala 64:55]
  assign _GEN_1025 = 11'h401 == fractionSum[12:2] ? 10'h200 : _GEN_1024; // @[Multiplier.scala 64:55]
  assign _GEN_1026 = 11'h402 == fractionSum[12:2] ? 10'h201 : _GEN_1025; // @[Multiplier.scala 64:55]
  assign _GEN_1027 = 11'h403 == fractionSum[12:2] ? 10'h201 : _GEN_1026; // @[Multiplier.scala 64:55]
  assign _GEN_1028 = 11'h404 == fractionSum[12:2] ? 10'h201 : _GEN_1027; // @[Multiplier.scala 64:55]
  assign _GEN_1029 = 11'h405 == fractionSum[12:2] ? 10'h202 : _GEN_1028; // @[Multiplier.scala 64:55]
  assign _GEN_1030 = 11'h406 == fractionSum[12:2] ? 10'h202 : _GEN_1029; // @[Multiplier.scala 64:55]
  assign _GEN_1031 = 11'h407 == fractionSum[12:2] ? 10'h202 : _GEN_1030; // @[Multiplier.scala 64:55]
  assign _GEN_1032 = 11'h408 == fractionSum[12:2] ? 10'h203 : _GEN_1031; // @[Multiplier.scala 64:55]
  assign _GEN_1033 = 11'h409 == fractionSum[12:2] ? 10'h203 : _GEN_1032; // @[Multiplier.scala 64:55]
  assign _GEN_1034 = 11'h40a == fractionSum[12:2] ? 10'h203 : _GEN_1033; // @[Multiplier.scala 64:55]
  assign _GEN_1035 = 11'h40b == fractionSum[12:2] ? 10'h204 : _GEN_1034; // @[Multiplier.scala 64:55]
  assign _GEN_1036 = 11'h40c == fractionSum[12:2] ? 10'h204 : _GEN_1035; // @[Multiplier.scala 64:55]
  assign _GEN_1037 = 11'h40d == fractionSum[12:2] ? 10'h205 : _GEN_1036; // @[Multiplier.scala 64:55]
  assign _GEN_1038 = 11'h40e == fractionSum[12:2] ? 10'h205 : _GEN_1037; // @[Multiplier.scala 64:55]
  assign _GEN_1039 = 11'h40f == fractionSum[12:2] ? 10'h205 : _GEN_1038; // @[Multiplier.scala 64:55]
  assign _GEN_1040 = 11'h410 == fractionSum[12:2] ? 10'h206 : _GEN_1039; // @[Multiplier.scala 64:55]
  assign _GEN_1041 = 11'h411 == fractionSum[12:2] ? 10'h206 : _GEN_1040; // @[Multiplier.scala 64:55]
  assign _GEN_1042 = 11'h412 == fractionSum[12:2] ? 10'h206 : _GEN_1041; // @[Multiplier.scala 64:55]
  assign _GEN_1043 = 11'h413 == fractionSum[12:2] ? 10'h207 : _GEN_1042; // @[Multiplier.scala 64:55]
  assign _GEN_1044 = 11'h414 == fractionSum[12:2] ? 10'h207 : _GEN_1043; // @[Multiplier.scala 64:55]
  assign _GEN_1045 = 11'h415 == fractionSum[12:2] ? 10'h207 : _GEN_1044; // @[Multiplier.scala 64:55]
  assign _GEN_1046 = 11'h416 == fractionSum[12:2] ? 10'h208 : _GEN_1045; // @[Multiplier.scala 64:55]
  assign _GEN_1047 = 11'h417 == fractionSum[12:2] ? 10'h208 : _GEN_1046; // @[Multiplier.scala 64:55]
  assign _GEN_1048 = 11'h418 == fractionSum[12:2] ? 10'h208 : _GEN_1047; // @[Multiplier.scala 64:55]
  assign _GEN_1049 = 11'h419 == fractionSum[12:2] ? 10'h209 : _GEN_1048; // @[Multiplier.scala 64:55]
  assign _GEN_1050 = 11'h41a == fractionSum[12:2] ? 10'h209 : _GEN_1049; // @[Multiplier.scala 64:55]
  assign _GEN_1051 = 11'h41b == fractionSum[12:2] ? 10'h209 : _GEN_1050; // @[Multiplier.scala 64:55]
  assign _GEN_1052 = 11'h41c == fractionSum[12:2] ? 10'h20a : _GEN_1051; // @[Multiplier.scala 64:55]
  assign _GEN_1053 = 11'h41d == fractionSum[12:2] ? 10'h20a : _GEN_1052; // @[Multiplier.scala 64:55]
  assign _GEN_1054 = 11'h41e == fractionSum[12:2] ? 10'h20b : _GEN_1053; // @[Multiplier.scala 64:55]
  assign _GEN_1055 = 11'h41f == fractionSum[12:2] ? 10'h20b : _GEN_1054; // @[Multiplier.scala 64:55]
  assign _GEN_1056 = 11'h420 == fractionSum[12:2] ? 10'h20b : _GEN_1055; // @[Multiplier.scala 64:55]
  assign _GEN_1057 = 11'h421 == fractionSum[12:2] ? 10'h20c : _GEN_1056; // @[Multiplier.scala 64:55]
  assign _GEN_1058 = 11'h422 == fractionSum[12:2] ? 10'h20c : _GEN_1057; // @[Multiplier.scala 64:55]
  assign _GEN_1059 = 11'h423 == fractionSum[12:2] ? 10'h20c : _GEN_1058; // @[Multiplier.scala 64:55]
  assign _GEN_1060 = 11'h424 == fractionSum[12:2] ? 10'h20d : _GEN_1059; // @[Multiplier.scala 64:55]
  assign _GEN_1061 = 11'h425 == fractionSum[12:2] ? 10'h20d : _GEN_1060; // @[Multiplier.scala 64:55]
  assign _GEN_1062 = 11'h426 == fractionSum[12:2] ? 10'h20d : _GEN_1061; // @[Multiplier.scala 64:55]
  assign _GEN_1063 = 11'h427 == fractionSum[12:2] ? 10'h20e : _GEN_1062; // @[Multiplier.scala 64:55]
  assign _GEN_1064 = 11'h428 == fractionSum[12:2] ? 10'h20e : _GEN_1063; // @[Multiplier.scala 64:55]
  assign _GEN_1065 = 11'h429 == fractionSum[12:2] ? 10'h20e : _GEN_1064; // @[Multiplier.scala 64:55]
  assign _GEN_1066 = 11'h42a == fractionSum[12:2] ? 10'h20f : _GEN_1065; // @[Multiplier.scala 64:55]
  assign _GEN_1067 = 11'h42b == fractionSum[12:2] ? 10'h20f : _GEN_1066; // @[Multiplier.scala 64:55]
  assign _GEN_1068 = 11'h42c == fractionSum[12:2] ? 10'h20f : _GEN_1067; // @[Multiplier.scala 64:55]
  assign _GEN_1069 = 11'h42d == fractionSum[12:2] ? 10'h210 : _GEN_1068; // @[Multiplier.scala 64:55]
  assign _GEN_1070 = 11'h42e == fractionSum[12:2] ? 10'h210 : _GEN_1069; // @[Multiplier.scala 64:55]
  assign _GEN_1071 = 11'h42f == fractionSum[12:2] ? 10'h211 : _GEN_1070; // @[Multiplier.scala 64:55]
  assign _GEN_1072 = 11'h430 == fractionSum[12:2] ? 10'h211 : _GEN_1071; // @[Multiplier.scala 64:55]
  assign _GEN_1073 = 11'h431 == fractionSum[12:2] ? 10'h211 : _GEN_1072; // @[Multiplier.scala 64:55]
  assign _GEN_1074 = 11'h432 == fractionSum[12:2] ? 10'h212 : _GEN_1073; // @[Multiplier.scala 64:55]
  assign _GEN_1075 = 11'h433 == fractionSum[12:2] ? 10'h212 : _GEN_1074; // @[Multiplier.scala 64:55]
  assign _GEN_1076 = 11'h434 == fractionSum[12:2] ? 10'h212 : _GEN_1075; // @[Multiplier.scala 64:55]
  assign _GEN_1077 = 11'h435 == fractionSum[12:2] ? 10'h213 : _GEN_1076; // @[Multiplier.scala 64:55]
  assign _GEN_1078 = 11'h436 == fractionSum[12:2] ? 10'h213 : _GEN_1077; // @[Multiplier.scala 64:55]
  assign _GEN_1079 = 11'h437 == fractionSum[12:2] ? 10'h213 : _GEN_1078; // @[Multiplier.scala 64:55]
  assign _GEN_1080 = 11'h438 == fractionSum[12:2] ? 10'h214 : _GEN_1079; // @[Multiplier.scala 64:55]
  assign _GEN_1081 = 11'h439 == fractionSum[12:2] ? 10'h214 : _GEN_1080; // @[Multiplier.scala 64:55]
  assign _GEN_1082 = 11'h43a == fractionSum[12:2] ? 10'h215 : _GEN_1081; // @[Multiplier.scala 64:55]
  assign _GEN_1083 = 11'h43b == fractionSum[12:2] ? 10'h215 : _GEN_1082; // @[Multiplier.scala 64:55]
  assign _GEN_1084 = 11'h43c == fractionSum[12:2] ? 10'h215 : _GEN_1083; // @[Multiplier.scala 64:55]
  assign _GEN_1085 = 11'h43d == fractionSum[12:2] ? 10'h216 : _GEN_1084; // @[Multiplier.scala 64:55]
  assign _GEN_1086 = 11'h43e == fractionSum[12:2] ? 10'h216 : _GEN_1085; // @[Multiplier.scala 64:55]
  assign _GEN_1087 = 11'h43f == fractionSum[12:2] ? 10'h216 : _GEN_1086; // @[Multiplier.scala 64:55]
  assign _GEN_1088 = 11'h440 == fractionSum[12:2] ? 10'h217 : _GEN_1087; // @[Multiplier.scala 64:55]
  assign _GEN_1089 = 11'h441 == fractionSum[12:2] ? 10'h217 : _GEN_1088; // @[Multiplier.scala 64:55]
  assign _GEN_1090 = 11'h442 == fractionSum[12:2] ? 10'h217 : _GEN_1089; // @[Multiplier.scala 64:55]
  assign _GEN_1091 = 11'h443 == fractionSum[12:2] ? 10'h218 : _GEN_1090; // @[Multiplier.scala 64:55]
  assign _GEN_1092 = 11'h444 == fractionSum[12:2] ? 10'h218 : _GEN_1091; // @[Multiplier.scala 64:55]
  assign _GEN_1093 = 11'h445 == fractionSum[12:2] ? 10'h218 : _GEN_1092; // @[Multiplier.scala 64:55]
  assign _GEN_1094 = 11'h446 == fractionSum[12:2] ? 10'h219 : _GEN_1093; // @[Multiplier.scala 64:55]
  assign _GEN_1095 = 11'h447 == fractionSum[12:2] ? 10'h219 : _GEN_1094; // @[Multiplier.scala 64:55]
  assign _GEN_1096 = 11'h448 == fractionSum[12:2] ? 10'h21a : _GEN_1095; // @[Multiplier.scala 64:55]
  assign _GEN_1097 = 11'h449 == fractionSum[12:2] ? 10'h21a : _GEN_1096; // @[Multiplier.scala 64:55]
  assign _GEN_1098 = 11'h44a == fractionSum[12:2] ? 10'h21a : _GEN_1097; // @[Multiplier.scala 64:55]
  assign _GEN_1099 = 11'h44b == fractionSum[12:2] ? 10'h21b : _GEN_1098; // @[Multiplier.scala 64:55]
  assign _GEN_1100 = 11'h44c == fractionSum[12:2] ? 10'h21b : _GEN_1099; // @[Multiplier.scala 64:55]
  assign _GEN_1101 = 11'h44d == fractionSum[12:2] ? 10'h21b : _GEN_1100; // @[Multiplier.scala 64:55]
  assign _GEN_1102 = 11'h44e == fractionSum[12:2] ? 10'h21c : _GEN_1101; // @[Multiplier.scala 64:55]
  assign _GEN_1103 = 11'h44f == fractionSum[12:2] ? 10'h21c : _GEN_1102; // @[Multiplier.scala 64:55]
  assign _GEN_1104 = 11'h450 == fractionSum[12:2] ? 10'h21c : _GEN_1103; // @[Multiplier.scala 64:55]
  assign _GEN_1105 = 11'h451 == fractionSum[12:2] ? 10'h21d : _GEN_1104; // @[Multiplier.scala 64:55]
  assign _GEN_1106 = 11'h452 == fractionSum[12:2] ? 10'h21d : _GEN_1105; // @[Multiplier.scala 64:55]
  assign _GEN_1107 = 11'h453 == fractionSum[12:2] ? 10'h21e : _GEN_1106; // @[Multiplier.scala 64:55]
  assign _GEN_1108 = 11'h454 == fractionSum[12:2] ? 10'h21e : _GEN_1107; // @[Multiplier.scala 64:55]
  assign _GEN_1109 = 11'h455 == fractionSum[12:2] ? 10'h21e : _GEN_1108; // @[Multiplier.scala 64:55]
  assign _GEN_1110 = 11'h456 == fractionSum[12:2] ? 10'h21f : _GEN_1109; // @[Multiplier.scala 64:55]
  assign _GEN_1111 = 11'h457 == fractionSum[12:2] ? 10'h21f : _GEN_1110; // @[Multiplier.scala 64:55]
  assign _GEN_1112 = 11'h458 == fractionSum[12:2] ? 10'h21f : _GEN_1111; // @[Multiplier.scala 64:55]
  assign _GEN_1113 = 11'h459 == fractionSum[12:2] ? 10'h220 : _GEN_1112; // @[Multiplier.scala 64:55]
  assign _GEN_1114 = 11'h45a == fractionSum[12:2] ? 10'h220 : _GEN_1113; // @[Multiplier.scala 64:55]
  assign _GEN_1115 = 11'h45b == fractionSum[12:2] ? 10'h221 : _GEN_1114; // @[Multiplier.scala 64:55]
  assign _GEN_1116 = 11'h45c == fractionSum[12:2] ? 10'h221 : _GEN_1115; // @[Multiplier.scala 64:55]
  assign _GEN_1117 = 11'h45d == fractionSum[12:2] ? 10'h221 : _GEN_1116; // @[Multiplier.scala 64:55]
  assign _GEN_1118 = 11'h45e == fractionSum[12:2] ? 10'h222 : _GEN_1117; // @[Multiplier.scala 64:55]
  assign _GEN_1119 = 11'h45f == fractionSum[12:2] ? 10'h222 : _GEN_1118; // @[Multiplier.scala 64:55]
  assign _GEN_1120 = 11'h460 == fractionSum[12:2] ? 10'h222 : _GEN_1119; // @[Multiplier.scala 64:55]
  assign _GEN_1121 = 11'h461 == fractionSum[12:2] ? 10'h223 : _GEN_1120; // @[Multiplier.scala 64:55]
  assign _GEN_1122 = 11'h462 == fractionSum[12:2] ? 10'h223 : _GEN_1121; // @[Multiplier.scala 64:55]
  assign _GEN_1123 = 11'h463 == fractionSum[12:2] ? 10'h223 : _GEN_1122; // @[Multiplier.scala 64:55]
  assign _GEN_1124 = 11'h464 == fractionSum[12:2] ? 10'h224 : _GEN_1123; // @[Multiplier.scala 64:55]
  assign _GEN_1125 = 11'h465 == fractionSum[12:2] ? 10'h224 : _GEN_1124; // @[Multiplier.scala 64:55]
  assign _GEN_1126 = 11'h466 == fractionSum[12:2] ? 10'h225 : _GEN_1125; // @[Multiplier.scala 64:55]
  assign _GEN_1127 = 11'h467 == fractionSum[12:2] ? 10'h225 : _GEN_1126; // @[Multiplier.scala 64:55]
  assign _GEN_1128 = 11'h468 == fractionSum[12:2] ? 10'h225 : _GEN_1127; // @[Multiplier.scala 64:55]
  assign _GEN_1129 = 11'h469 == fractionSum[12:2] ? 10'h226 : _GEN_1128; // @[Multiplier.scala 64:55]
  assign _GEN_1130 = 11'h46a == fractionSum[12:2] ? 10'h226 : _GEN_1129; // @[Multiplier.scala 64:55]
  assign _GEN_1131 = 11'h46b == fractionSum[12:2] ? 10'h226 : _GEN_1130; // @[Multiplier.scala 64:55]
  assign _GEN_1132 = 11'h46c == fractionSum[12:2] ? 10'h227 : _GEN_1131; // @[Multiplier.scala 64:55]
  assign _GEN_1133 = 11'h46d == fractionSum[12:2] ? 10'h227 : _GEN_1132; // @[Multiplier.scala 64:55]
  assign _GEN_1134 = 11'h46e == fractionSum[12:2] ? 10'h228 : _GEN_1133; // @[Multiplier.scala 64:55]
  assign _GEN_1135 = 11'h46f == fractionSum[12:2] ? 10'h228 : _GEN_1134; // @[Multiplier.scala 64:55]
  assign _GEN_1136 = 11'h470 == fractionSum[12:2] ? 10'h228 : _GEN_1135; // @[Multiplier.scala 64:55]
  assign _GEN_1137 = 11'h471 == fractionSum[12:2] ? 10'h229 : _GEN_1136; // @[Multiplier.scala 64:55]
  assign _GEN_1138 = 11'h472 == fractionSum[12:2] ? 10'h229 : _GEN_1137; // @[Multiplier.scala 64:55]
  assign _GEN_1139 = 11'h473 == fractionSum[12:2] ? 10'h229 : _GEN_1138; // @[Multiplier.scala 64:55]
  assign _GEN_1140 = 11'h474 == fractionSum[12:2] ? 10'h22a : _GEN_1139; // @[Multiplier.scala 64:55]
  assign _GEN_1141 = 11'h475 == fractionSum[12:2] ? 10'h22a : _GEN_1140; // @[Multiplier.scala 64:55]
  assign _GEN_1142 = 11'h476 == fractionSum[12:2] ? 10'h22b : _GEN_1141; // @[Multiplier.scala 64:55]
  assign _GEN_1143 = 11'h477 == fractionSum[12:2] ? 10'h22b : _GEN_1142; // @[Multiplier.scala 64:55]
  assign _GEN_1144 = 11'h478 == fractionSum[12:2] ? 10'h22b : _GEN_1143; // @[Multiplier.scala 64:55]
  assign _GEN_1145 = 11'h479 == fractionSum[12:2] ? 10'h22c : _GEN_1144; // @[Multiplier.scala 64:55]
  assign _GEN_1146 = 11'h47a == fractionSum[12:2] ? 10'h22c : _GEN_1145; // @[Multiplier.scala 64:55]
  assign _GEN_1147 = 11'h47b == fractionSum[12:2] ? 10'h22c : _GEN_1146; // @[Multiplier.scala 64:55]
  assign _GEN_1148 = 11'h47c == fractionSum[12:2] ? 10'h22d : _GEN_1147; // @[Multiplier.scala 64:55]
  assign _GEN_1149 = 11'h47d == fractionSum[12:2] ? 10'h22d : _GEN_1148; // @[Multiplier.scala 64:55]
  assign _GEN_1150 = 11'h47e == fractionSum[12:2] ? 10'h22e : _GEN_1149; // @[Multiplier.scala 64:55]
  assign _GEN_1151 = 11'h47f == fractionSum[12:2] ? 10'h22e : _GEN_1150; // @[Multiplier.scala 64:55]
  assign _GEN_1152 = 11'h480 == fractionSum[12:2] ? 10'h22e : _GEN_1151; // @[Multiplier.scala 64:55]
  assign _GEN_1153 = 11'h481 == fractionSum[12:2] ? 10'h22f : _GEN_1152; // @[Multiplier.scala 64:55]
  assign _GEN_1154 = 11'h482 == fractionSum[12:2] ? 10'h22f : _GEN_1153; // @[Multiplier.scala 64:55]
  assign _GEN_1155 = 11'h483 == fractionSum[12:2] ? 10'h22f : _GEN_1154; // @[Multiplier.scala 64:55]
  assign _GEN_1156 = 11'h484 == fractionSum[12:2] ? 10'h230 : _GEN_1155; // @[Multiplier.scala 64:55]
  assign _GEN_1157 = 11'h485 == fractionSum[12:2] ? 10'h230 : _GEN_1156; // @[Multiplier.scala 64:55]
  assign _GEN_1158 = 11'h486 == fractionSum[12:2] ? 10'h231 : _GEN_1157; // @[Multiplier.scala 64:55]
  assign _GEN_1159 = 11'h487 == fractionSum[12:2] ? 10'h231 : _GEN_1158; // @[Multiplier.scala 64:55]
  assign _GEN_1160 = 11'h488 == fractionSum[12:2] ? 10'h231 : _GEN_1159; // @[Multiplier.scala 64:55]
  assign _GEN_1161 = 11'h489 == fractionSum[12:2] ? 10'h232 : _GEN_1160; // @[Multiplier.scala 64:55]
  assign _GEN_1162 = 11'h48a == fractionSum[12:2] ? 10'h232 : _GEN_1161; // @[Multiplier.scala 64:55]
  assign _GEN_1163 = 11'h48b == fractionSum[12:2] ? 10'h233 : _GEN_1162; // @[Multiplier.scala 64:55]
  assign _GEN_1164 = 11'h48c == fractionSum[12:2] ? 10'h233 : _GEN_1163; // @[Multiplier.scala 64:55]
  assign _GEN_1165 = 11'h48d == fractionSum[12:2] ? 10'h233 : _GEN_1164; // @[Multiplier.scala 64:55]
  assign _GEN_1166 = 11'h48e == fractionSum[12:2] ? 10'h234 : _GEN_1165; // @[Multiplier.scala 64:55]
  assign _GEN_1167 = 11'h48f == fractionSum[12:2] ? 10'h234 : _GEN_1166; // @[Multiplier.scala 64:55]
  assign _GEN_1168 = 11'h490 == fractionSum[12:2] ? 10'h234 : _GEN_1167; // @[Multiplier.scala 64:55]
  assign _GEN_1169 = 11'h491 == fractionSum[12:2] ? 10'h235 : _GEN_1168; // @[Multiplier.scala 64:55]
  assign _GEN_1170 = 11'h492 == fractionSum[12:2] ? 10'h235 : _GEN_1169; // @[Multiplier.scala 64:55]
  assign _GEN_1171 = 11'h493 == fractionSum[12:2] ? 10'h236 : _GEN_1170; // @[Multiplier.scala 64:55]
  assign _GEN_1172 = 11'h494 == fractionSum[12:2] ? 10'h236 : _GEN_1171; // @[Multiplier.scala 64:55]
  assign _GEN_1173 = 11'h495 == fractionSum[12:2] ? 10'h236 : _GEN_1172; // @[Multiplier.scala 64:55]
  assign _GEN_1174 = 11'h496 == fractionSum[12:2] ? 10'h237 : _GEN_1173; // @[Multiplier.scala 64:55]
  assign _GEN_1175 = 11'h497 == fractionSum[12:2] ? 10'h237 : _GEN_1174; // @[Multiplier.scala 64:55]
  assign _GEN_1176 = 11'h498 == fractionSum[12:2] ? 10'h237 : _GEN_1175; // @[Multiplier.scala 64:55]
  assign _GEN_1177 = 11'h499 == fractionSum[12:2] ? 10'h238 : _GEN_1176; // @[Multiplier.scala 64:55]
  assign _GEN_1178 = 11'h49a == fractionSum[12:2] ? 10'h238 : _GEN_1177; // @[Multiplier.scala 64:55]
  assign _GEN_1179 = 11'h49b == fractionSum[12:2] ? 10'h239 : _GEN_1178; // @[Multiplier.scala 64:55]
  assign _GEN_1180 = 11'h49c == fractionSum[12:2] ? 10'h239 : _GEN_1179; // @[Multiplier.scala 64:55]
  assign _GEN_1181 = 11'h49d == fractionSum[12:2] ? 10'h239 : _GEN_1180; // @[Multiplier.scala 64:55]
  assign _GEN_1182 = 11'h49e == fractionSum[12:2] ? 10'h23a : _GEN_1181; // @[Multiplier.scala 64:55]
  assign _GEN_1183 = 11'h49f == fractionSum[12:2] ? 10'h23a : _GEN_1182; // @[Multiplier.scala 64:55]
  assign _GEN_1184 = 11'h4a0 == fractionSum[12:2] ? 10'h23b : _GEN_1183; // @[Multiplier.scala 64:55]
  assign _GEN_1185 = 11'h4a1 == fractionSum[12:2] ? 10'h23b : _GEN_1184; // @[Multiplier.scala 64:55]
  assign _GEN_1186 = 11'h4a2 == fractionSum[12:2] ? 10'h23b : _GEN_1185; // @[Multiplier.scala 64:55]
  assign _GEN_1187 = 11'h4a3 == fractionSum[12:2] ? 10'h23c : _GEN_1186; // @[Multiplier.scala 64:55]
  assign _GEN_1188 = 11'h4a4 == fractionSum[12:2] ? 10'h23c : _GEN_1187; // @[Multiplier.scala 64:55]
  assign _GEN_1189 = 11'h4a5 == fractionSum[12:2] ? 10'h23d : _GEN_1188; // @[Multiplier.scala 64:55]
  assign _GEN_1190 = 11'h4a6 == fractionSum[12:2] ? 10'h23d : _GEN_1189; // @[Multiplier.scala 64:55]
  assign _GEN_1191 = 11'h4a7 == fractionSum[12:2] ? 10'h23d : _GEN_1190; // @[Multiplier.scala 64:55]
  assign _GEN_1192 = 11'h4a8 == fractionSum[12:2] ? 10'h23e : _GEN_1191; // @[Multiplier.scala 64:55]
  assign _GEN_1193 = 11'h4a9 == fractionSum[12:2] ? 10'h23e : _GEN_1192; // @[Multiplier.scala 64:55]
  assign _GEN_1194 = 11'h4aa == fractionSum[12:2] ? 10'h23e : _GEN_1193; // @[Multiplier.scala 64:55]
  assign _GEN_1195 = 11'h4ab == fractionSum[12:2] ? 10'h23f : _GEN_1194; // @[Multiplier.scala 64:55]
  assign _GEN_1196 = 11'h4ac == fractionSum[12:2] ? 10'h23f : _GEN_1195; // @[Multiplier.scala 64:55]
  assign _GEN_1197 = 11'h4ad == fractionSum[12:2] ? 10'h240 : _GEN_1196; // @[Multiplier.scala 64:55]
  assign _GEN_1198 = 11'h4ae == fractionSum[12:2] ? 10'h240 : _GEN_1197; // @[Multiplier.scala 64:55]
  assign _GEN_1199 = 11'h4af == fractionSum[12:2] ? 10'h240 : _GEN_1198; // @[Multiplier.scala 64:55]
  assign _GEN_1200 = 11'h4b0 == fractionSum[12:2] ? 10'h241 : _GEN_1199; // @[Multiplier.scala 64:55]
  assign _GEN_1201 = 11'h4b1 == fractionSum[12:2] ? 10'h241 : _GEN_1200; // @[Multiplier.scala 64:55]
  assign _GEN_1202 = 11'h4b2 == fractionSum[12:2] ? 10'h242 : _GEN_1201; // @[Multiplier.scala 64:55]
  assign _GEN_1203 = 11'h4b3 == fractionSum[12:2] ? 10'h242 : _GEN_1202; // @[Multiplier.scala 64:55]
  assign _GEN_1204 = 11'h4b4 == fractionSum[12:2] ? 10'h242 : _GEN_1203; // @[Multiplier.scala 64:55]
  assign _GEN_1205 = 11'h4b5 == fractionSum[12:2] ? 10'h243 : _GEN_1204; // @[Multiplier.scala 64:55]
  assign _GEN_1206 = 11'h4b6 == fractionSum[12:2] ? 10'h243 : _GEN_1205; // @[Multiplier.scala 64:55]
  assign _GEN_1207 = 11'h4b7 == fractionSum[12:2] ? 10'h244 : _GEN_1206; // @[Multiplier.scala 64:55]
  assign _GEN_1208 = 11'h4b8 == fractionSum[12:2] ? 10'h244 : _GEN_1207; // @[Multiplier.scala 64:55]
  assign _GEN_1209 = 11'h4b9 == fractionSum[12:2] ? 10'h244 : _GEN_1208; // @[Multiplier.scala 64:55]
  assign _GEN_1210 = 11'h4ba == fractionSum[12:2] ? 10'h245 : _GEN_1209; // @[Multiplier.scala 64:55]
  assign _GEN_1211 = 11'h4bb == fractionSum[12:2] ? 10'h245 : _GEN_1210; // @[Multiplier.scala 64:55]
  assign _GEN_1212 = 11'h4bc == fractionSum[12:2] ? 10'h245 : _GEN_1211; // @[Multiplier.scala 64:55]
  assign _GEN_1213 = 11'h4bd == fractionSum[12:2] ? 10'h246 : _GEN_1212; // @[Multiplier.scala 64:55]
  assign _GEN_1214 = 11'h4be == fractionSum[12:2] ? 10'h246 : _GEN_1213; // @[Multiplier.scala 64:55]
  assign _GEN_1215 = 11'h4bf == fractionSum[12:2] ? 10'h247 : _GEN_1214; // @[Multiplier.scala 64:55]
  assign _GEN_1216 = 11'h4c0 == fractionSum[12:2] ? 10'h247 : _GEN_1215; // @[Multiplier.scala 64:55]
  assign _GEN_1217 = 11'h4c1 == fractionSum[12:2] ? 10'h247 : _GEN_1216; // @[Multiplier.scala 64:55]
  assign _GEN_1218 = 11'h4c2 == fractionSum[12:2] ? 10'h248 : _GEN_1217; // @[Multiplier.scala 64:55]
  assign _GEN_1219 = 11'h4c3 == fractionSum[12:2] ? 10'h248 : _GEN_1218; // @[Multiplier.scala 64:55]
  assign _GEN_1220 = 11'h4c4 == fractionSum[12:2] ? 10'h249 : _GEN_1219; // @[Multiplier.scala 64:55]
  assign _GEN_1221 = 11'h4c5 == fractionSum[12:2] ? 10'h249 : _GEN_1220; // @[Multiplier.scala 64:55]
  assign _GEN_1222 = 11'h4c6 == fractionSum[12:2] ? 10'h249 : _GEN_1221; // @[Multiplier.scala 64:55]
  assign _GEN_1223 = 11'h4c7 == fractionSum[12:2] ? 10'h24a : _GEN_1222; // @[Multiplier.scala 64:55]
  assign _GEN_1224 = 11'h4c8 == fractionSum[12:2] ? 10'h24a : _GEN_1223; // @[Multiplier.scala 64:55]
  assign _GEN_1225 = 11'h4c9 == fractionSum[12:2] ? 10'h24b : _GEN_1224; // @[Multiplier.scala 64:55]
  assign _GEN_1226 = 11'h4ca == fractionSum[12:2] ? 10'h24b : _GEN_1225; // @[Multiplier.scala 64:55]
  assign _GEN_1227 = 11'h4cb == fractionSum[12:2] ? 10'h24b : _GEN_1226; // @[Multiplier.scala 64:55]
  assign _GEN_1228 = 11'h4cc == fractionSum[12:2] ? 10'h24c : _GEN_1227; // @[Multiplier.scala 64:55]
  assign _GEN_1229 = 11'h4cd == fractionSum[12:2] ? 10'h24c : _GEN_1228; // @[Multiplier.scala 64:55]
  assign _GEN_1230 = 11'h4ce == fractionSum[12:2] ? 10'h24d : _GEN_1229; // @[Multiplier.scala 64:55]
  assign _GEN_1231 = 11'h4cf == fractionSum[12:2] ? 10'h24d : _GEN_1230; // @[Multiplier.scala 64:55]
  assign _GEN_1232 = 11'h4d0 == fractionSum[12:2] ? 10'h24d : _GEN_1231; // @[Multiplier.scala 64:55]
  assign _GEN_1233 = 11'h4d1 == fractionSum[12:2] ? 10'h24e : _GEN_1232; // @[Multiplier.scala 64:55]
  assign _GEN_1234 = 11'h4d2 == fractionSum[12:2] ? 10'h24e : _GEN_1233; // @[Multiplier.scala 64:55]
  assign _GEN_1235 = 11'h4d3 == fractionSum[12:2] ? 10'h24f : _GEN_1234; // @[Multiplier.scala 64:55]
  assign _GEN_1236 = 11'h4d4 == fractionSum[12:2] ? 10'h24f : _GEN_1235; // @[Multiplier.scala 64:55]
  assign _GEN_1237 = 11'h4d5 == fractionSum[12:2] ? 10'h24f : _GEN_1236; // @[Multiplier.scala 64:55]
  assign _GEN_1238 = 11'h4d6 == fractionSum[12:2] ? 10'h250 : _GEN_1237; // @[Multiplier.scala 64:55]
  assign _GEN_1239 = 11'h4d7 == fractionSum[12:2] ? 10'h250 : _GEN_1238; // @[Multiplier.scala 64:55]
  assign _GEN_1240 = 11'h4d8 == fractionSum[12:2] ? 10'h251 : _GEN_1239; // @[Multiplier.scala 64:55]
  assign _GEN_1241 = 11'h4d9 == fractionSum[12:2] ? 10'h251 : _GEN_1240; // @[Multiplier.scala 64:55]
  assign _GEN_1242 = 11'h4da == fractionSum[12:2] ? 10'h251 : _GEN_1241; // @[Multiplier.scala 64:55]
  assign _GEN_1243 = 11'h4db == fractionSum[12:2] ? 10'h252 : _GEN_1242; // @[Multiplier.scala 64:55]
  assign _GEN_1244 = 11'h4dc == fractionSum[12:2] ? 10'h252 : _GEN_1243; // @[Multiplier.scala 64:55]
  assign _GEN_1245 = 11'h4dd == fractionSum[12:2] ? 10'h253 : _GEN_1244; // @[Multiplier.scala 64:55]
  assign _GEN_1246 = 11'h4de == fractionSum[12:2] ? 10'h253 : _GEN_1245; // @[Multiplier.scala 64:55]
  assign _GEN_1247 = 11'h4df == fractionSum[12:2] ? 10'h253 : _GEN_1246; // @[Multiplier.scala 64:55]
  assign _GEN_1248 = 11'h4e0 == fractionSum[12:2] ? 10'h254 : _GEN_1247; // @[Multiplier.scala 64:55]
  assign _GEN_1249 = 11'h4e1 == fractionSum[12:2] ? 10'h254 : _GEN_1248; // @[Multiplier.scala 64:55]
  assign _GEN_1250 = 11'h4e2 == fractionSum[12:2] ? 10'h255 : _GEN_1249; // @[Multiplier.scala 64:55]
  assign _GEN_1251 = 11'h4e3 == fractionSum[12:2] ? 10'h255 : _GEN_1250; // @[Multiplier.scala 64:55]
  assign _GEN_1252 = 11'h4e4 == fractionSum[12:2] ? 10'h255 : _GEN_1251; // @[Multiplier.scala 64:55]
  assign _GEN_1253 = 11'h4e5 == fractionSum[12:2] ? 10'h256 : _GEN_1252; // @[Multiplier.scala 64:55]
  assign _GEN_1254 = 11'h4e6 == fractionSum[12:2] ? 10'h256 : _GEN_1253; // @[Multiplier.scala 64:55]
  assign _GEN_1255 = 11'h4e7 == fractionSum[12:2] ? 10'h257 : _GEN_1254; // @[Multiplier.scala 64:55]
  assign _GEN_1256 = 11'h4e8 == fractionSum[12:2] ? 10'h257 : _GEN_1255; // @[Multiplier.scala 64:55]
  assign _GEN_1257 = 11'h4e9 == fractionSum[12:2] ? 10'h257 : _GEN_1256; // @[Multiplier.scala 64:55]
  assign _GEN_1258 = 11'h4ea == fractionSum[12:2] ? 10'h258 : _GEN_1257; // @[Multiplier.scala 64:55]
  assign _GEN_1259 = 11'h4eb == fractionSum[12:2] ? 10'h258 : _GEN_1258; // @[Multiplier.scala 64:55]
  assign _GEN_1260 = 11'h4ec == fractionSum[12:2] ? 10'h259 : _GEN_1259; // @[Multiplier.scala 64:55]
  assign _GEN_1261 = 11'h4ed == fractionSum[12:2] ? 10'h259 : _GEN_1260; // @[Multiplier.scala 64:55]
  assign _GEN_1262 = 11'h4ee == fractionSum[12:2] ? 10'h25a : _GEN_1261; // @[Multiplier.scala 64:55]
  assign _GEN_1263 = 11'h4ef == fractionSum[12:2] ? 10'h25a : _GEN_1262; // @[Multiplier.scala 64:55]
  assign _GEN_1264 = 11'h4f0 == fractionSum[12:2] ? 10'h25a : _GEN_1263; // @[Multiplier.scala 64:55]
  assign _GEN_1265 = 11'h4f1 == fractionSum[12:2] ? 10'h25b : _GEN_1264; // @[Multiplier.scala 64:55]
  assign _GEN_1266 = 11'h4f2 == fractionSum[12:2] ? 10'h25b : _GEN_1265; // @[Multiplier.scala 64:55]
  assign _GEN_1267 = 11'h4f3 == fractionSum[12:2] ? 10'h25c : _GEN_1266; // @[Multiplier.scala 64:55]
  assign _GEN_1268 = 11'h4f4 == fractionSum[12:2] ? 10'h25c : _GEN_1267; // @[Multiplier.scala 64:55]
  assign _GEN_1269 = 11'h4f5 == fractionSum[12:2] ? 10'h25c : _GEN_1268; // @[Multiplier.scala 64:55]
  assign _GEN_1270 = 11'h4f6 == fractionSum[12:2] ? 10'h25d : _GEN_1269; // @[Multiplier.scala 64:55]
  assign _GEN_1271 = 11'h4f7 == fractionSum[12:2] ? 10'h25d : _GEN_1270; // @[Multiplier.scala 64:55]
  assign _GEN_1272 = 11'h4f8 == fractionSum[12:2] ? 10'h25e : _GEN_1271; // @[Multiplier.scala 64:55]
  assign _GEN_1273 = 11'h4f9 == fractionSum[12:2] ? 10'h25e : _GEN_1272; // @[Multiplier.scala 64:55]
  assign _GEN_1274 = 11'h4fa == fractionSum[12:2] ? 10'h25e : _GEN_1273; // @[Multiplier.scala 64:55]
  assign _GEN_1275 = 11'h4fb == fractionSum[12:2] ? 10'h25f : _GEN_1274; // @[Multiplier.scala 64:55]
  assign _GEN_1276 = 11'h4fc == fractionSum[12:2] ? 10'h25f : _GEN_1275; // @[Multiplier.scala 64:55]
  assign _GEN_1277 = 11'h4fd == fractionSum[12:2] ? 10'h260 : _GEN_1276; // @[Multiplier.scala 64:55]
  assign _GEN_1278 = 11'h4fe == fractionSum[12:2] ? 10'h260 : _GEN_1277; // @[Multiplier.scala 64:55]
  assign _GEN_1279 = 11'h4ff == fractionSum[12:2] ? 10'h260 : _GEN_1278; // @[Multiplier.scala 64:55]
  assign _GEN_1280 = 11'h500 == fractionSum[12:2] ? 10'h261 : _GEN_1279; // @[Multiplier.scala 64:55]
  assign _GEN_1281 = 11'h501 == fractionSum[12:2] ? 10'h261 : _GEN_1280; // @[Multiplier.scala 64:55]
  assign _GEN_1282 = 11'h502 == fractionSum[12:2] ? 10'h262 : _GEN_1281; // @[Multiplier.scala 64:55]
  assign _GEN_1283 = 11'h503 == fractionSum[12:2] ? 10'h262 : _GEN_1282; // @[Multiplier.scala 64:55]
  assign _GEN_1284 = 11'h504 == fractionSum[12:2] ? 10'h263 : _GEN_1283; // @[Multiplier.scala 64:55]
  assign _GEN_1285 = 11'h505 == fractionSum[12:2] ? 10'h263 : _GEN_1284; // @[Multiplier.scala 64:55]
  assign _GEN_1286 = 11'h506 == fractionSum[12:2] ? 10'h263 : _GEN_1285; // @[Multiplier.scala 64:55]
  assign _GEN_1287 = 11'h507 == fractionSum[12:2] ? 10'h264 : _GEN_1286; // @[Multiplier.scala 64:55]
  assign _GEN_1288 = 11'h508 == fractionSum[12:2] ? 10'h264 : _GEN_1287; // @[Multiplier.scala 64:55]
  assign _GEN_1289 = 11'h509 == fractionSum[12:2] ? 10'h265 : _GEN_1288; // @[Multiplier.scala 64:55]
  assign _GEN_1290 = 11'h50a == fractionSum[12:2] ? 10'h265 : _GEN_1289; // @[Multiplier.scala 64:55]
  assign _GEN_1291 = 11'h50b == fractionSum[12:2] ? 10'h265 : _GEN_1290; // @[Multiplier.scala 64:55]
  assign _GEN_1292 = 11'h50c == fractionSum[12:2] ? 10'h266 : _GEN_1291; // @[Multiplier.scala 64:55]
  assign _GEN_1293 = 11'h50d == fractionSum[12:2] ? 10'h266 : _GEN_1292; // @[Multiplier.scala 64:55]
  assign _GEN_1294 = 11'h50e == fractionSum[12:2] ? 10'h267 : _GEN_1293; // @[Multiplier.scala 64:55]
  assign _GEN_1295 = 11'h50f == fractionSum[12:2] ? 10'h267 : _GEN_1294; // @[Multiplier.scala 64:55]
  assign _GEN_1296 = 11'h510 == fractionSum[12:2] ? 10'h268 : _GEN_1295; // @[Multiplier.scala 64:55]
  assign _GEN_1297 = 11'h511 == fractionSum[12:2] ? 10'h268 : _GEN_1296; // @[Multiplier.scala 64:55]
  assign _GEN_1298 = 11'h512 == fractionSum[12:2] ? 10'h268 : _GEN_1297; // @[Multiplier.scala 64:55]
  assign _GEN_1299 = 11'h513 == fractionSum[12:2] ? 10'h269 : _GEN_1298; // @[Multiplier.scala 64:55]
  assign _GEN_1300 = 11'h514 == fractionSum[12:2] ? 10'h269 : _GEN_1299; // @[Multiplier.scala 64:55]
  assign _GEN_1301 = 11'h515 == fractionSum[12:2] ? 10'h26a : _GEN_1300; // @[Multiplier.scala 64:55]
  assign _GEN_1302 = 11'h516 == fractionSum[12:2] ? 10'h26a : _GEN_1301; // @[Multiplier.scala 64:55]
  assign _GEN_1303 = 11'h517 == fractionSum[12:2] ? 10'h26a : _GEN_1302; // @[Multiplier.scala 64:55]
  assign _GEN_1304 = 11'h518 == fractionSum[12:2] ? 10'h26b : _GEN_1303; // @[Multiplier.scala 64:55]
  assign _GEN_1305 = 11'h519 == fractionSum[12:2] ? 10'h26b : _GEN_1304; // @[Multiplier.scala 64:55]
  assign _GEN_1306 = 11'h51a == fractionSum[12:2] ? 10'h26c : _GEN_1305; // @[Multiplier.scala 64:55]
  assign _GEN_1307 = 11'h51b == fractionSum[12:2] ? 10'h26c : _GEN_1306; // @[Multiplier.scala 64:55]
  assign _GEN_1308 = 11'h51c == fractionSum[12:2] ? 10'h26d : _GEN_1307; // @[Multiplier.scala 64:55]
  assign _GEN_1309 = 11'h51d == fractionSum[12:2] ? 10'h26d : _GEN_1308; // @[Multiplier.scala 64:55]
  assign _GEN_1310 = 11'h51e == fractionSum[12:2] ? 10'h26d : _GEN_1309; // @[Multiplier.scala 64:55]
  assign _GEN_1311 = 11'h51f == fractionSum[12:2] ? 10'h26e : _GEN_1310; // @[Multiplier.scala 64:55]
  assign _GEN_1312 = 11'h520 == fractionSum[12:2] ? 10'h26e : _GEN_1311; // @[Multiplier.scala 64:55]
  assign _GEN_1313 = 11'h521 == fractionSum[12:2] ? 10'h26f : _GEN_1312; // @[Multiplier.scala 64:55]
  assign _GEN_1314 = 11'h522 == fractionSum[12:2] ? 10'h26f : _GEN_1313; // @[Multiplier.scala 64:55]
  assign _GEN_1315 = 11'h523 == fractionSum[12:2] ? 10'h26f : _GEN_1314; // @[Multiplier.scala 64:55]
  assign _GEN_1316 = 11'h524 == fractionSum[12:2] ? 10'h270 : _GEN_1315; // @[Multiplier.scala 64:55]
  assign _GEN_1317 = 11'h525 == fractionSum[12:2] ? 10'h270 : _GEN_1316; // @[Multiplier.scala 64:55]
  assign _GEN_1318 = 11'h526 == fractionSum[12:2] ? 10'h271 : _GEN_1317; // @[Multiplier.scala 64:55]
  assign _GEN_1319 = 11'h527 == fractionSum[12:2] ? 10'h271 : _GEN_1318; // @[Multiplier.scala 64:55]
  assign _GEN_1320 = 11'h528 == fractionSum[12:2] ? 10'h272 : _GEN_1319; // @[Multiplier.scala 64:55]
  assign _GEN_1321 = 11'h529 == fractionSum[12:2] ? 10'h272 : _GEN_1320; // @[Multiplier.scala 64:55]
  assign _GEN_1322 = 11'h52a == fractionSum[12:2] ? 10'h272 : _GEN_1321; // @[Multiplier.scala 64:55]
  assign _GEN_1323 = 11'h52b == fractionSum[12:2] ? 10'h273 : _GEN_1322; // @[Multiplier.scala 64:55]
  assign _GEN_1324 = 11'h52c == fractionSum[12:2] ? 10'h273 : _GEN_1323; // @[Multiplier.scala 64:55]
  assign _GEN_1325 = 11'h52d == fractionSum[12:2] ? 10'h274 : _GEN_1324; // @[Multiplier.scala 64:55]
  assign _GEN_1326 = 11'h52e == fractionSum[12:2] ? 10'h274 : _GEN_1325; // @[Multiplier.scala 64:55]
  assign _GEN_1327 = 11'h52f == fractionSum[12:2] ? 10'h275 : _GEN_1326; // @[Multiplier.scala 64:55]
  assign _GEN_1328 = 11'h530 == fractionSum[12:2] ? 10'h275 : _GEN_1327; // @[Multiplier.scala 64:55]
  assign _GEN_1329 = 11'h531 == fractionSum[12:2] ? 10'h275 : _GEN_1328; // @[Multiplier.scala 64:55]
  assign _GEN_1330 = 11'h532 == fractionSum[12:2] ? 10'h276 : _GEN_1329; // @[Multiplier.scala 64:55]
  assign _GEN_1331 = 11'h533 == fractionSum[12:2] ? 10'h276 : _GEN_1330; // @[Multiplier.scala 64:55]
  assign _GEN_1332 = 11'h534 == fractionSum[12:2] ? 10'h277 : _GEN_1331; // @[Multiplier.scala 64:55]
  assign _GEN_1333 = 11'h535 == fractionSum[12:2] ? 10'h277 : _GEN_1332; // @[Multiplier.scala 64:55]
  assign _GEN_1334 = 11'h536 == fractionSum[12:2] ? 10'h278 : _GEN_1333; // @[Multiplier.scala 64:55]
  assign _GEN_1335 = 11'h537 == fractionSum[12:2] ? 10'h278 : _GEN_1334; // @[Multiplier.scala 64:55]
  assign _GEN_1336 = 11'h538 == fractionSum[12:2] ? 10'h278 : _GEN_1335; // @[Multiplier.scala 64:55]
  assign _GEN_1337 = 11'h539 == fractionSum[12:2] ? 10'h279 : _GEN_1336; // @[Multiplier.scala 64:55]
  assign _GEN_1338 = 11'h53a == fractionSum[12:2] ? 10'h279 : _GEN_1337; // @[Multiplier.scala 64:55]
  assign _GEN_1339 = 11'h53b == fractionSum[12:2] ? 10'h27a : _GEN_1338; // @[Multiplier.scala 64:55]
  assign _GEN_1340 = 11'h53c == fractionSum[12:2] ? 10'h27a : _GEN_1339; // @[Multiplier.scala 64:55]
  assign _GEN_1341 = 11'h53d == fractionSum[12:2] ? 10'h27b : _GEN_1340; // @[Multiplier.scala 64:55]
  assign _GEN_1342 = 11'h53e == fractionSum[12:2] ? 10'h27b : _GEN_1341; // @[Multiplier.scala 64:55]
  assign _GEN_1343 = 11'h53f == fractionSum[12:2] ? 10'h27b : _GEN_1342; // @[Multiplier.scala 64:55]
  assign _GEN_1344 = 11'h540 == fractionSum[12:2] ? 10'h27c : _GEN_1343; // @[Multiplier.scala 64:55]
  assign _GEN_1345 = 11'h541 == fractionSum[12:2] ? 10'h27c : _GEN_1344; // @[Multiplier.scala 64:55]
  assign _GEN_1346 = 11'h542 == fractionSum[12:2] ? 10'h27d : _GEN_1345; // @[Multiplier.scala 64:55]
  assign _GEN_1347 = 11'h543 == fractionSum[12:2] ? 10'h27d : _GEN_1346; // @[Multiplier.scala 64:55]
  assign _GEN_1348 = 11'h544 == fractionSum[12:2] ? 10'h27e : _GEN_1347; // @[Multiplier.scala 64:55]
  assign _GEN_1349 = 11'h545 == fractionSum[12:2] ? 10'h27e : _GEN_1348; // @[Multiplier.scala 64:55]
  assign _GEN_1350 = 11'h546 == fractionSum[12:2] ? 10'h27e : _GEN_1349; // @[Multiplier.scala 64:55]
  assign _GEN_1351 = 11'h547 == fractionSum[12:2] ? 10'h27f : _GEN_1350; // @[Multiplier.scala 64:55]
  assign _GEN_1352 = 11'h548 == fractionSum[12:2] ? 10'h27f : _GEN_1351; // @[Multiplier.scala 64:55]
  assign _GEN_1353 = 11'h549 == fractionSum[12:2] ? 10'h280 : _GEN_1352; // @[Multiplier.scala 64:55]
  assign _GEN_1354 = 11'h54a == fractionSum[12:2] ? 10'h280 : _GEN_1353; // @[Multiplier.scala 64:55]
  assign _GEN_1355 = 11'h54b == fractionSum[12:2] ? 10'h281 : _GEN_1354; // @[Multiplier.scala 64:55]
  assign _GEN_1356 = 11'h54c == fractionSum[12:2] ? 10'h281 : _GEN_1355; // @[Multiplier.scala 64:55]
  assign _GEN_1357 = 11'h54d == fractionSum[12:2] ? 10'h281 : _GEN_1356; // @[Multiplier.scala 64:55]
  assign _GEN_1358 = 11'h54e == fractionSum[12:2] ? 10'h282 : _GEN_1357; // @[Multiplier.scala 64:55]
  assign _GEN_1359 = 11'h54f == fractionSum[12:2] ? 10'h282 : _GEN_1358; // @[Multiplier.scala 64:55]
  assign _GEN_1360 = 11'h550 == fractionSum[12:2] ? 10'h283 : _GEN_1359; // @[Multiplier.scala 64:55]
  assign _GEN_1361 = 11'h551 == fractionSum[12:2] ? 10'h283 : _GEN_1360; // @[Multiplier.scala 64:55]
  assign _GEN_1362 = 11'h552 == fractionSum[12:2] ? 10'h284 : _GEN_1361; // @[Multiplier.scala 64:55]
  assign _GEN_1363 = 11'h553 == fractionSum[12:2] ? 10'h284 : _GEN_1362; // @[Multiplier.scala 64:55]
  assign _GEN_1364 = 11'h554 == fractionSum[12:2] ? 10'h284 : _GEN_1363; // @[Multiplier.scala 64:55]
  assign _GEN_1365 = 11'h555 == fractionSum[12:2] ? 10'h285 : _GEN_1364; // @[Multiplier.scala 64:55]
  assign _GEN_1366 = 11'h556 == fractionSum[12:2] ? 10'h285 : _GEN_1365; // @[Multiplier.scala 64:55]
  assign _GEN_1367 = 11'h557 == fractionSum[12:2] ? 10'h286 : _GEN_1366; // @[Multiplier.scala 64:55]
  assign _GEN_1368 = 11'h558 == fractionSum[12:2] ? 10'h286 : _GEN_1367; // @[Multiplier.scala 64:55]
  assign _GEN_1369 = 11'h559 == fractionSum[12:2] ? 10'h287 : _GEN_1368; // @[Multiplier.scala 64:55]
  assign _GEN_1370 = 11'h55a == fractionSum[12:2] ? 10'h287 : _GEN_1369; // @[Multiplier.scala 64:55]
  assign _GEN_1371 = 11'h55b == fractionSum[12:2] ? 10'h288 : _GEN_1370; // @[Multiplier.scala 64:55]
  assign _GEN_1372 = 11'h55c == fractionSum[12:2] ? 10'h288 : _GEN_1371; // @[Multiplier.scala 64:55]
  assign _GEN_1373 = 11'h55d == fractionSum[12:2] ? 10'h288 : _GEN_1372; // @[Multiplier.scala 64:55]
  assign _GEN_1374 = 11'h55e == fractionSum[12:2] ? 10'h289 : _GEN_1373; // @[Multiplier.scala 64:55]
  assign _GEN_1375 = 11'h55f == fractionSum[12:2] ? 10'h289 : _GEN_1374; // @[Multiplier.scala 64:55]
  assign _GEN_1376 = 11'h560 == fractionSum[12:2] ? 10'h28a : _GEN_1375; // @[Multiplier.scala 64:55]
  assign _GEN_1377 = 11'h561 == fractionSum[12:2] ? 10'h28a : _GEN_1376; // @[Multiplier.scala 64:55]
  assign _GEN_1378 = 11'h562 == fractionSum[12:2] ? 10'h28b : _GEN_1377; // @[Multiplier.scala 64:55]
  assign _GEN_1379 = 11'h563 == fractionSum[12:2] ? 10'h28b : _GEN_1378; // @[Multiplier.scala 64:55]
  assign _GEN_1380 = 11'h564 == fractionSum[12:2] ? 10'h28c : _GEN_1379; // @[Multiplier.scala 64:55]
  assign _GEN_1381 = 11'h565 == fractionSum[12:2] ? 10'h28c : _GEN_1380; // @[Multiplier.scala 64:55]
  assign _GEN_1382 = 11'h566 == fractionSum[12:2] ? 10'h28c : _GEN_1381; // @[Multiplier.scala 64:55]
  assign _GEN_1383 = 11'h567 == fractionSum[12:2] ? 10'h28d : _GEN_1382; // @[Multiplier.scala 64:55]
  assign _GEN_1384 = 11'h568 == fractionSum[12:2] ? 10'h28d : _GEN_1383; // @[Multiplier.scala 64:55]
  assign _GEN_1385 = 11'h569 == fractionSum[12:2] ? 10'h28e : _GEN_1384; // @[Multiplier.scala 64:55]
  assign _GEN_1386 = 11'h56a == fractionSum[12:2] ? 10'h28e : _GEN_1385; // @[Multiplier.scala 64:55]
  assign _GEN_1387 = 11'h56b == fractionSum[12:2] ? 10'h28f : _GEN_1386; // @[Multiplier.scala 64:55]
  assign _GEN_1388 = 11'h56c == fractionSum[12:2] ? 10'h28f : _GEN_1387; // @[Multiplier.scala 64:55]
  assign _GEN_1389 = 11'h56d == fractionSum[12:2] ? 10'h28f : _GEN_1388; // @[Multiplier.scala 64:55]
  assign _GEN_1390 = 11'h56e == fractionSum[12:2] ? 10'h290 : _GEN_1389; // @[Multiplier.scala 64:55]
  assign _GEN_1391 = 11'h56f == fractionSum[12:2] ? 10'h290 : _GEN_1390; // @[Multiplier.scala 64:55]
  assign _GEN_1392 = 11'h570 == fractionSum[12:2] ? 10'h291 : _GEN_1391; // @[Multiplier.scala 64:55]
  assign _GEN_1393 = 11'h571 == fractionSum[12:2] ? 10'h291 : _GEN_1392; // @[Multiplier.scala 64:55]
  assign _GEN_1394 = 11'h572 == fractionSum[12:2] ? 10'h292 : _GEN_1393; // @[Multiplier.scala 64:55]
  assign _GEN_1395 = 11'h573 == fractionSum[12:2] ? 10'h292 : _GEN_1394; // @[Multiplier.scala 64:55]
  assign _GEN_1396 = 11'h574 == fractionSum[12:2] ? 10'h293 : _GEN_1395; // @[Multiplier.scala 64:55]
  assign _GEN_1397 = 11'h575 == fractionSum[12:2] ? 10'h293 : _GEN_1396; // @[Multiplier.scala 64:55]
  assign _GEN_1398 = 11'h576 == fractionSum[12:2] ? 10'h294 : _GEN_1397; // @[Multiplier.scala 64:55]
  assign _GEN_1399 = 11'h577 == fractionSum[12:2] ? 10'h294 : _GEN_1398; // @[Multiplier.scala 64:55]
  assign _GEN_1400 = 11'h578 == fractionSum[12:2] ? 10'h294 : _GEN_1399; // @[Multiplier.scala 64:55]
  assign _GEN_1401 = 11'h579 == fractionSum[12:2] ? 10'h295 : _GEN_1400; // @[Multiplier.scala 64:55]
  assign _GEN_1402 = 11'h57a == fractionSum[12:2] ? 10'h295 : _GEN_1401; // @[Multiplier.scala 64:55]
  assign _GEN_1403 = 11'h57b == fractionSum[12:2] ? 10'h296 : _GEN_1402; // @[Multiplier.scala 64:55]
  assign _GEN_1404 = 11'h57c == fractionSum[12:2] ? 10'h296 : _GEN_1403; // @[Multiplier.scala 64:55]
  assign _GEN_1405 = 11'h57d == fractionSum[12:2] ? 10'h297 : _GEN_1404; // @[Multiplier.scala 64:55]
  assign _GEN_1406 = 11'h57e == fractionSum[12:2] ? 10'h297 : _GEN_1405; // @[Multiplier.scala 64:55]
  assign _GEN_1407 = 11'h57f == fractionSum[12:2] ? 10'h298 : _GEN_1406; // @[Multiplier.scala 64:55]
  assign _GEN_1408 = 11'h580 == fractionSum[12:2] ? 10'h298 : _GEN_1407; // @[Multiplier.scala 64:55]
  assign _GEN_1409 = 11'h581 == fractionSum[12:2] ? 10'h298 : _GEN_1408; // @[Multiplier.scala 64:55]
  assign _GEN_1410 = 11'h582 == fractionSum[12:2] ? 10'h299 : _GEN_1409; // @[Multiplier.scala 64:55]
  assign _GEN_1411 = 11'h583 == fractionSum[12:2] ? 10'h299 : _GEN_1410; // @[Multiplier.scala 64:55]
  assign _GEN_1412 = 11'h584 == fractionSum[12:2] ? 10'h29a : _GEN_1411; // @[Multiplier.scala 64:55]
  assign _GEN_1413 = 11'h585 == fractionSum[12:2] ? 10'h29a : _GEN_1412; // @[Multiplier.scala 64:55]
  assign _GEN_1414 = 11'h586 == fractionSum[12:2] ? 10'h29b : _GEN_1413; // @[Multiplier.scala 64:55]
  assign _GEN_1415 = 11'h587 == fractionSum[12:2] ? 10'h29b : _GEN_1414; // @[Multiplier.scala 64:55]
  assign _GEN_1416 = 11'h588 == fractionSum[12:2] ? 10'h29c : _GEN_1415; // @[Multiplier.scala 64:55]
  assign _GEN_1417 = 11'h589 == fractionSum[12:2] ? 10'h29c : _GEN_1416; // @[Multiplier.scala 64:55]
  assign _GEN_1418 = 11'h58a == fractionSum[12:2] ? 10'h29c : _GEN_1417; // @[Multiplier.scala 64:55]
  assign _GEN_1419 = 11'h58b == fractionSum[12:2] ? 10'h29d : _GEN_1418; // @[Multiplier.scala 64:55]
  assign _GEN_1420 = 11'h58c == fractionSum[12:2] ? 10'h29d : _GEN_1419; // @[Multiplier.scala 64:55]
  assign _GEN_1421 = 11'h58d == fractionSum[12:2] ? 10'h29e : _GEN_1420; // @[Multiplier.scala 64:55]
  assign _GEN_1422 = 11'h58e == fractionSum[12:2] ? 10'h29e : _GEN_1421; // @[Multiplier.scala 64:55]
  assign _GEN_1423 = 11'h58f == fractionSum[12:2] ? 10'h29f : _GEN_1422; // @[Multiplier.scala 64:55]
  assign _GEN_1424 = 11'h590 == fractionSum[12:2] ? 10'h29f : _GEN_1423; // @[Multiplier.scala 64:55]
  assign _GEN_1425 = 11'h591 == fractionSum[12:2] ? 10'h2a0 : _GEN_1424; // @[Multiplier.scala 64:55]
  assign _GEN_1426 = 11'h592 == fractionSum[12:2] ? 10'h2a0 : _GEN_1425; // @[Multiplier.scala 64:55]
  assign _GEN_1427 = 11'h593 == fractionSum[12:2] ? 10'h2a1 : _GEN_1426; // @[Multiplier.scala 64:55]
  assign _GEN_1428 = 11'h594 == fractionSum[12:2] ? 10'h2a1 : _GEN_1427; // @[Multiplier.scala 64:55]
  assign _GEN_1429 = 11'h595 == fractionSum[12:2] ? 10'h2a1 : _GEN_1428; // @[Multiplier.scala 64:55]
  assign _GEN_1430 = 11'h596 == fractionSum[12:2] ? 10'h2a2 : _GEN_1429; // @[Multiplier.scala 64:55]
  assign _GEN_1431 = 11'h597 == fractionSum[12:2] ? 10'h2a2 : _GEN_1430; // @[Multiplier.scala 64:55]
  assign _GEN_1432 = 11'h598 == fractionSum[12:2] ? 10'h2a3 : _GEN_1431; // @[Multiplier.scala 64:55]
  assign _GEN_1433 = 11'h599 == fractionSum[12:2] ? 10'h2a3 : _GEN_1432; // @[Multiplier.scala 64:55]
  assign _GEN_1434 = 11'h59a == fractionSum[12:2] ? 10'h2a4 : _GEN_1433; // @[Multiplier.scala 64:55]
  assign _GEN_1435 = 11'h59b == fractionSum[12:2] ? 10'h2a4 : _GEN_1434; // @[Multiplier.scala 64:55]
  assign _GEN_1436 = 11'h59c == fractionSum[12:2] ? 10'h2a5 : _GEN_1435; // @[Multiplier.scala 64:55]
  assign _GEN_1437 = 11'h59d == fractionSum[12:2] ? 10'h2a5 : _GEN_1436; // @[Multiplier.scala 64:55]
  assign _GEN_1438 = 11'h59e == fractionSum[12:2] ? 10'h2a6 : _GEN_1437; // @[Multiplier.scala 64:55]
  assign _GEN_1439 = 11'h59f == fractionSum[12:2] ? 10'h2a6 : _GEN_1438; // @[Multiplier.scala 64:55]
  assign _GEN_1440 = 11'h5a0 == fractionSum[12:2] ? 10'h2a7 : _GEN_1439; // @[Multiplier.scala 64:55]
  assign _GEN_1441 = 11'h5a1 == fractionSum[12:2] ? 10'h2a7 : _GEN_1440; // @[Multiplier.scala 64:55]
  assign _GEN_1442 = 11'h5a2 == fractionSum[12:2] ? 10'h2a7 : _GEN_1441; // @[Multiplier.scala 64:55]
  assign _GEN_1443 = 11'h5a3 == fractionSum[12:2] ? 10'h2a8 : _GEN_1442; // @[Multiplier.scala 64:55]
  assign _GEN_1444 = 11'h5a4 == fractionSum[12:2] ? 10'h2a8 : _GEN_1443; // @[Multiplier.scala 64:55]
  assign _GEN_1445 = 11'h5a5 == fractionSum[12:2] ? 10'h2a9 : _GEN_1444; // @[Multiplier.scala 64:55]
  assign _GEN_1446 = 11'h5a6 == fractionSum[12:2] ? 10'h2a9 : _GEN_1445; // @[Multiplier.scala 64:55]
  assign _GEN_1447 = 11'h5a7 == fractionSum[12:2] ? 10'h2aa : _GEN_1446; // @[Multiplier.scala 64:55]
  assign _GEN_1448 = 11'h5a8 == fractionSum[12:2] ? 10'h2aa : _GEN_1447; // @[Multiplier.scala 64:55]
  assign _GEN_1449 = 11'h5a9 == fractionSum[12:2] ? 10'h2ab : _GEN_1448; // @[Multiplier.scala 64:55]
  assign _GEN_1450 = 11'h5aa == fractionSum[12:2] ? 10'h2ab : _GEN_1449; // @[Multiplier.scala 64:55]
  assign _GEN_1451 = 11'h5ab == fractionSum[12:2] ? 10'h2ac : _GEN_1450; // @[Multiplier.scala 64:55]
  assign _GEN_1452 = 11'h5ac == fractionSum[12:2] ? 10'h2ac : _GEN_1451; // @[Multiplier.scala 64:55]
  assign _GEN_1453 = 11'h5ad == fractionSum[12:2] ? 10'h2ad : _GEN_1452; // @[Multiplier.scala 64:55]
  assign _GEN_1454 = 11'h5ae == fractionSum[12:2] ? 10'h2ad : _GEN_1453; // @[Multiplier.scala 64:55]
  assign _GEN_1455 = 11'h5af == fractionSum[12:2] ? 10'h2ad : _GEN_1454; // @[Multiplier.scala 64:55]
  assign _GEN_1456 = 11'h5b0 == fractionSum[12:2] ? 10'h2ae : _GEN_1455; // @[Multiplier.scala 64:55]
  assign _GEN_1457 = 11'h5b1 == fractionSum[12:2] ? 10'h2ae : _GEN_1456; // @[Multiplier.scala 64:55]
  assign _GEN_1458 = 11'h5b2 == fractionSum[12:2] ? 10'h2af : _GEN_1457; // @[Multiplier.scala 64:55]
  assign _GEN_1459 = 11'h5b3 == fractionSum[12:2] ? 10'h2af : _GEN_1458; // @[Multiplier.scala 64:55]
  assign _GEN_1460 = 11'h5b4 == fractionSum[12:2] ? 10'h2b0 : _GEN_1459; // @[Multiplier.scala 64:55]
  assign _GEN_1461 = 11'h5b5 == fractionSum[12:2] ? 10'h2b0 : _GEN_1460; // @[Multiplier.scala 64:55]
  assign _GEN_1462 = 11'h5b6 == fractionSum[12:2] ? 10'h2b1 : _GEN_1461; // @[Multiplier.scala 64:55]
  assign _GEN_1463 = 11'h5b7 == fractionSum[12:2] ? 10'h2b1 : _GEN_1462; // @[Multiplier.scala 64:55]
  assign _GEN_1464 = 11'h5b8 == fractionSum[12:2] ? 10'h2b2 : _GEN_1463; // @[Multiplier.scala 64:55]
  assign _GEN_1465 = 11'h5b9 == fractionSum[12:2] ? 10'h2b2 : _GEN_1464; // @[Multiplier.scala 64:55]
  assign _GEN_1466 = 11'h5ba == fractionSum[12:2] ? 10'h2b3 : _GEN_1465; // @[Multiplier.scala 64:55]
  assign _GEN_1467 = 11'h5bb == fractionSum[12:2] ? 10'h2b3 : _GEN_1466; // @[Multiplier.scala 64:55]
  assign _GEN_1468 = 11'h5bc == fractionSum[12:2] ? 10'h2b4 : _GEN_1467; // @[Multiplier.scala 64:55]
  assign _GEN_1469 = 11'h5bd == fractionSum[12:2] ? 10'h2b4 : _GEN_1468; // @[Multiplier.scala 64:55]
  assign _GEN_1470 = 11'h5be == fractionSum[12:2] ? 10'h2b4 : _GEN_1469; // @[Multiplier.scala 64:55]
  assign _GEN_1471 = 11'h5bf == fractionSum[12:2] ? 10'h2b5 : _GEN_1470; // @[Multiplier.scala 64:55]
  assign _GEN_1472 = 11'h5c0 == fractionSum[12:2] ? 10'h2b5 : _GEN_1471; // @[Multiplier.scala 64:55]
  assign _GEN_1473 = 11'h5c1 == fractionSum[12:2] ? 10'h2b6 : _GEN_1472; // @[Multiplier.scala 64:55]
  assign _GEN_1474 = 11'h5c2 == fractionSum[12:2] ? 10'h2b6 : _GEN_1473; // @[Multiplier.scala 64:55]
  assign _GEN_1475 = 11'h5c3 == fractionSum[12:2] ? 10'h2b7 : _GEN_1474; // @[Multiplier.scala 64:55]
  assign _GEN_1476 = 11'h5c4 == fractionSum[12:2] ? 10'h2b7 : _GEN_1475; // @[Multiplier.scala 64:55]
  assign _GEN_1477 = 11'h5c5 == fractionSum[12:2] ? 10'h2b8 : _GEN_1476; // @[Multiplier.scala 64:55]
  assign _GEN_1478 = 11'h5c6 == fractionSum[12:2] ? 10'h2b8 : _GEN_1477; // @[Multiplier.scala 64:55]
  assign _GEN_1479 = 11'h5c7 == fractionSum[12:2] ? 10'h2b9 : _GEN_1478; // @[Multiplier.scala 64:55]
  assign _GEN_1480 = 11'h5c8 == fractionSum[12:2] ? 10'h2b9 : _GEN_1479; // @[Multiplier.scala 64:55]
  assign _GEN_1481 = 11'h5c9 == fractionSum[12:2] ? 10'h2ba : _GEN_1480; // @[Multiplier.scala 64:55]
  assign _GEN_1482 = 11'h5ca == fractionSum[12:2] ? 10'h2ba : _GEN_1481; // @[Multiplier.scala 64:55]
  assign _GEN_1483 = 11'h5cb == fractionSum[12:2] ? 10'h2bb : _GEN_1482; // @[Multiplier.scala 64:55]
  assign _GEN_1484 = 11'h5cc == fractionSum[12:2] ? 10'h2bb : _GEN_1483; // @[Multiplier.scala 64:55]
  assign _GEN_1485 = 11'h5cd == fractionSum[12:2] ? 10'h2bc : _GEN_1484; // @[Multiplier.scala 64:55]
  assign _GEN_1486 = 11'h5ce == fractionSum[12:2] ? 10'h2bc : _GEN_1485; // @[Multiplier.scala 64:55]
  assign _GEN_1487 = 11'h5cf == fractionSum[12:2] ? 10'h2bc : _GEN_1486; // @[Multiplier.scala 64:55]
  assign _GEN_1488 = 11'h5d0 == fractionSum[12:2] ? 10'h2bd : _GEN_1487; // @[Multiplier.scala 64:55]
  assign _GEN_1489 = 11'h5d1 == fractionSum[12:2] ? 10'h2bd : _GEN_1488; // @[Multiplier.scala 64:55]
  assign _GEN_1490 = 11'h5d2 == fractionSum[12:2] ? 10'h2be : _GEN_1489; // @[Multiplier.scala 64:55]
  assign _GEN_1491 = 11'h5d3 == fractionSum[12:2] ? 10'h2be : _GEN_1490; // @[Multiplier.scala 64:55]
  assign _GEN_1492 = 11'h5d4 == fractionSum[12:2] ? 10'h2bf : _GEN_1491; // @[Multiplier.scala 64:55]
  assign _GEN_1493 = 11'h5d5 == fractionSum[12:2] ? 10'h2bf : _GEN_1492; // @[Multiplier.scala 64:55]
  assign _GEN_1494 = 11'h5d6 == fractionSum[12:2] ? 10'h2c0 : _GEN_1493; // @[Multiplier.scala 64:55]
  assign _GEN_1495 = 11'h5d7 == fractionSum[12:2] ? 10'h2c0 : _GEN_1494; // @[Multiplier.scala 64:55]
  assign _GEN_1496 = 11'h5d8 == fractionSum[12:2] ? 10'h2c1 : _GEN_1495; // @[Multiplier.scala 64:55]
  assign _GEN_1497 = 11'h5d9 == fractionSum[12:2] ? 10'h2c1 : _GEN_1496; // @[Multiplier.scala 64:55]
  assign _GEN_1498 = 11'h5da == fractionSum[12:2] ? 10'h2c2 : _GEN_1497; // @[Multiplier.scala 64:55]
  assign _GEN_1499 = 11'h5db == fractionSum[12:2] ? 10'h2c2 : _GEN_1498; // @[Multiplier.scala 64:55]
  assign _GEN_1500 = 11'h5dc == fractionSum[12:2] ? 10'h2c3 : _GEN_1499; // @[Multiplier.scala 64:55]
  assign _GEN_1501 = 11'h5dd == fractionSum[12:2] ? 10'h2c3 : _GEN_1500; // @[Multiplier.scala 64:55]
  assign _GEN_1502 = 11'h5de == fractionSum[12:2] ? 10'h2c4 : _GEN_1501; // @[Multiplier.scala 64:55]
  assign _GEN_1503 = 11'h5df == fractionSum[12:2] ? 10'h2c4 : _GEN_1502; // @[Multiplier.scala 64:55]
  assign _GEN_1504 = 11'h5e0 == fractionSum[12:2] ? 10'h2c5 : _GEN_1503; // @[Multiplier.scala 64:55]
  assign _GEN_1505 = 11'h5e1 == fractionSum[12:2] ? 10'h2c5 : _GEN_1504; // @[Multiplier.scala 64:55]
  assign _GEN_1506 = 11'h5e2 == fractionSum[12:2] ? 10'h2c6 : _GEN_1505; // @[Multiplier.scala 64:55]
  assign _GEN_1507 = 11'h5e3 == fractionSum[12:2] ? 10'h2c6 : _GEN_1506; // @[Multiplier.scala 64:55]
  assign _GEN_1508 = 11'h5e4 == fractionSum[12:2] ? 10'h2c6 : _GEN_1507; // @[Multiplier.scala 64:55]
  assign _GEN_1509 = 11'h5e5 == fractionSum[12:2] ? 10'h2c7 : _GEN_1508; // @[Multiplier.scala 64:55]
  assign _GEN_1510 = 11'h5e6 == fractionSum[12:2] ? 10'h2c7 : _GEN_1509; // @[Multiplier.scala 64:55]
  assign _GEN_1511 = 11'h5e7 == fractionSum[12:2] ? 10'h2c8 : _GEN_1510; // @[Multiplier.scala 64:55]
  assign _GEN_1512 = 11'h5e8 == fractionSum[12:2] ? 10'h2c8 : _GEN_1511; // @[Multiplier.scala 64:55]
  assign _GEN_1513 = 11'h5e9 == fractionSum[12:2] ? 10'h2c9 : _GEN_1512; // @[Multiplier.scala 64:55]
  assign _GEN_1514 = 11'h5ea == fractionSum[12:2] ? 10'h2c9 : _GEN_1513; // @[Multiplier.scala 64:55]
  assign _GEN_1515 = 11'h5eb == fractionSum[12:2] ? 10'h2ca : _GEN_1514; // @[Multiplier.scala 64:55]
  assign _GEN_1516 = 11'h5ec == fractionSum[12:2] ? 10'h2ca : _GEN_1515; // @[Multiplier.scala 64:55]
  assign _GEN_1517 = 11'h5ed == fractionSum[12:2] ? 10'h2cb : _GEN_1516; // @[Multiplier.scala 64:55]
  assign _GEN_1518 = 11'h5ee == fractionSum[12:2] ? 10'h2cb : _GEN_1517; // @[Multiplier.scala 64:55]
  assign _GEN_1519 = 11'h5ef == fractionSum[12:2] ? 10'h2cc : _GEN_1518; // @[Multiplier.scala 64:55]
  assign _GEN_1520 = 11'h5f0 == fractionSum[12:2] ? 10'h2cc : _GEN_1519; // @[Multiplier.scala 64:55]
  assign _GEN_1521 = 11'h5f1 == fractionSum[12:2] ? 10'h2cd : _GEN_1520; // @[Multiplier.scala 64:55]
  assign _GEN_1522 = 11'h5f2 == fractionSum[12:2] ? 10'h2cd : _GEN_1521; // @[Multiplier.scala 64:55]
  assign _GEN_1523 = 11'h5f3 == fractionSum[12:2] ? 10'h2ce : _GEN_1522; // @[Multiplier.scala 64:55]
  assign _GEN_1524 = 11'h5f4 == fractionSum[12:2] ? 10'h2ce : _GEN_1523; // @[Multiplier.scala 64:55]
  assign _GEN_1525 = 11'h5f5 == fractionSum[12:2] ? 10'h2cf : _GEN_1524; // @[Multiplier.scala 64:55]
  assign _GEN_1526 = 11'h5f6 == fractionSum[12:2] ? 10'h2cf : _GEN_1525; // @[Multiplier.scala 64:55]
  assign _GEN_1527 = 11'h5f7 == fractionSum[12:2] ? 10'h2d0 : _GEN_1526; // @[Multiplier.scala 64:55]
  assign _GEN_1528 = 11'h5f8 == fractionSum[12:2] ? 10'h2d0 : _GEN_1527; // @[Multiplier.scala 64:55]
  assign _GEN_1529 = 11'h5f9 == fractionSum[12:2] ? 10'h2d1 : _GEN_1528; // @[Multiplier.scala 64:55]
  assign _GEN_1530 = 11'h5fa == fractionSum[12:2] ? 10'h2d1 : _GEN_1529; // @[Multiplier.scala 64:55]
  assign _GEN_1531 = 11'h5fb == fractionSum[12:2] ? 10'h2d2 : _GEN_1530; // @[Multiplier.scala 64:55]
  assign _GEN_1532 = 11'h5fc == fractionSum[12:2] ? 10'h2d2 : _GEN_1531; // @[Multiplier.scala 64:55]
  assign _GEN_1533 = 11'h5fd == fractionSum[12:2] ? 10'h2d3 : _GEN_1532; // @[Multiplier.scala 64:55]
  assign _GEN_1534 = 11'h5fe == fractionSum[12:2] ? 10'h2d3 : _GEN_1533; // @[Multiplier.scala 64:55]
  assign _GEN_1535 = 11'h5ff == fractionSum[12:2] ? 10'h2d4 : _GEN_1534; // @[Multiplier.scala 64:55]
  assign _GEN_1536 = 11'h600 == fractionSum[12:2] ? 10'h2d4 : _GEN_1535; // @[Multiplier.scala 64:55]
  assign _GEN_1537 = 11'h601 == fractionSum[12:2] ? 10'h2d5 : _GEN_1536; // @[Multiplier.scala 64:55]
  assign _GEN_1538 = 11'h602 == fractionSum[12:2] ? 10'h2d5 : _GEN_1537; // @[Multiplier.scala 64:55]
  assign _GEN_1539 = 11'h603 == fractionSum[12:2] ? 10'h2d6 : _GEN_1538; // @[Multiplier.scala 64:55]
  assign _GEN_1540 = 11'h604 == fractionSum[12:2] ? 10'h2d6 : _GEN_1539; // @[Multiplier.scala 64:55]
  assign _GEN_1541 = 11'h605 == fractionSum[12:2] ? 10'h2d7 : _GEN_1540; // @[Multiplier.scala 64:55]
  assign _GEN_1542 = 11'h606 == fractionSum[12:2] ? 10'h2d7 : _GEN_1541; // @[Multiplier.scala 64:55]
  assign _GEN_1543 = 11'h607 == fractionSum[12:2] ? 10'h2d8 : _GEN_1542; // @[Multiplier.scala 64:55]
  assign _GEN_1544 = 11'h608 == fractionSum[12:2] ? 10'h2d8 : _GEN_1543; // @[Multiplier.scala 64:55]
  assign _GEN_1545 = 11'h609 == fractionSum[12:2] ? 10'h2d9 : _GEN_1544; // @[Multiplier.scala 64:55]
  assign _GEN_1546 = 11'h60a == fractionSum[12:2] ? 10'h2d9 : _GEN_1545; // @[Multiplier.scala 64:55]
  assign _GEN_1547 = 11'h60b == fractionSum[12:2] ? 10'h2d9 : _GEN_1546; // @[Multiplier.scala 64:55]
  assign _GEN_1548 = 11'h60c == fractionSum[12:2] ? 10'h2da : _GEN_1547; // @[Multiplier.scala 64:55]
  assign _GEN_1549 = 11'h60d == fractionSum[12:2] ? 10'h2da : _GEN_1548; // @[Multiplier.scala 64:55]
  assign _GEN_1550 = 11'h60e == fractionSum[12:2] ? 10'h2db : _GEN_1549; // @[Multiplier.scala 64:55]
  assign _GEN_1551 = 11'h60f == fractionSum[12:2] ? 10'h2db : _GEN_1550; // @[Multiplier.scala 64:55]
  assign _GEN_1552 = 11'h610 == fractionSum[12:2] ? 10'h2dc : _GEN_1551; // @[Multiplier.scala 64:55]
  assign _GEN_1553 = 11'h611 == fractionSum[12:2] ? 10'h2dc : _GEN_1552; // @[Multiplier.scala 64:55]
  assign _GEN_1554 = 11'h612 == fractionSum[12:2] ? 10'h2dd : _GEN_1553; // @[Multiplier.scala 64:55]
  assign _GEN_1555 = 11'h613 == fractionSum[12:2] ? 10'h2dd : _GEN_1554; // @[Multiplier.scala 64:55]
  assign _GEN_1556 = 11'h614 == fractionSum[12:2] ? 10'h2de : _GEN_1555; // @[Multiplier.scala 64:55]
  assign _GEN_1557 = 11'h615 == fractionSum[12:2] ? 10'h2de : _GEN_1556; // @[Multiplier.scala 64:55]
  assign _GEN_1558 = 11'h616 == fractionSum[12:2] ? 10'h2df : _GEN_1557; // @[Multiplier.scala 64:55]
  assign _GEN_1559 = 11'h617 == fractionSum[12:2] ? 10'h2df : _GEN_1558; // @[Multiplier.scala 64:55]
  assign _GEN_1560 = 11'h618 == fractionSum[12:2] ? 10'h2e0 : _GEN_1559; // @[Multiplier.scala 64:55]
  assign _GEN_1561 = 11'h619 == fractionSum[12:2] ? 10'h2e0 : _GEN_1560; // @[Multiplier.scala 64:55]
  assign _GEN_1562 = 11'h61a == fractionSum[12:2] ? 10'h2e1 : _GEN_1561; // @[Multiplier.scala 64:55]
  assign _GEN_1563 = 11'h61b == fractionSum[12:2] ? 10'h2e1 : _GEN_1562; // @[Multiplier.scala 64:55]
  assign _GEN_1564 = 11'h61c == fractionSum[12:2] ? 10'h2e2 : _GEN_1563; // @[Multiplier.scala 64:55]
  assign _GEN_1565 = 11'h61d == fractionSum[12:2] ? 10'h2e2 : _GEN_1564; // @[Multiplier.scala 64:55]
  assign _GEN_1566 = 11'h61e == fractionSum[12:2] ? 10'h2e3 : _GEN_1565; // @[Multiplier.scala 64:55]
  assign _GEN_1567 = 11'h61f == fractionSum[12:2] ? 10'h2e3 : _GEN_1566; // @[Multiplier.scala 64:55]
  assign _GEN_1568 = 11'h620 == fractionSum[12:2] ? 10'h2e4 : _GEN_1567; // @[Multiplier.scala 64:55]
  assign _GEN_1569 = 11'h621 == fractionSum[12:2] ? 10'h2e4 : _GEN_1568; // @[Multiplier.scala 64:55]
  assign _GEN_1570 = 11'h622 == fractionSum[12:2] ? 10'h2e5 : _GEN_1569; // @[Multiplier.scala 64:55]
  assign _GEN_1571 = 11'h623 == fractionSum[12:2] ? 10'h2e5 : _GEN_1570; // @[Multiplier.scala 64:55]
  assign _GEN_1572 = 11'h624 == fractionSum[12:2] ? 10'h2e6 : _GEN_1571; // @[Multiplier.scala 64:55]
  assign _GEN_1573 = 11'h625 == fractionSum[12:2] ? 10'h2e6 : _GEN_1572; // @[Multiplier.scala 64:55]
  assign _GEN_1574 = 11'h626 == fractionSum[12:2] ? 10'h2e7 : _GEN_1573; // @[Multiplier.scala 64:55]
  assign _GEN_1575 = 11'h627 == fractionSum[12:2] ? 10'h2e7 : _GEN_1574; // @[Multiplier.scala 64:55]
  assign _GEN_1576 = 11'h628 == fractionSum[12:2] ? 10'h2e8 : _GEN_1575; // @[Multiplier.scala 64:55]
  assign _GEN_1577 = 11'h629 == fractionSum[12:2] ? 10'h2e8 : _GEN_1576; // @[Multiplier.scala 64:55]
  assign _GEN_1578 = 11'h62a == fractionSum[12:2] ? 10'h2e9 : _GEN_1577; // @[Multiplier.scala 64:55]
  assign _GEN_1579 = 11'h62b == fractionSum[12:2] ? 10'h2e9 : _GEN_1578; // @[Multiplier.scala 64:55]
  assign _GEN_1580 = 11'h62c == fractionSum[12:2] ? 10'h2ea : _GEN_1579; // @[Multiplier.scala 64:55]
  assign _GEN_1581 = 11'h62d == fractionSum[12:2] ? 10'h2ea : _GEN_1580; // @[Multiplier.scala 64:55]
  assign _GEN_1582 = 11'h62e == fractionSum[12:2] ? 10'h2eb : _GEN_1581; // @[Multiplier.scala 64:55]
  assign _GEN_1583 = 11'h62f == fractionSum[12:2] ? 10'h2eb : _GEN_1582; // @[Multiplier.scala 64:55]
  assign _GEN_1584 = 11'h630 == fractionSum[12:2] ? 10'h2ec : _GEN_1583; // @[Multiplier.scala 64:55]
  assign _GEN_1585 = 11'h631 == fractionSum[12:2] ? 10'h2ec : _GEN_1584; // @[Multiplier.scala 64:55]
  assign _GEN_1586 = 11'h632 == fractionSum[12:2] ? 10'h2ed : _GEN_1585; // @[Multiplier.scala 64:55]
  assign _GEN_1587 = 11'h633 == fractionSum[12:2] ? 10'h2ee : _GEN_1586; // @[Multiplier.scala 64:55]
  assign _GEN_1588 = 11'h634 == fractionSum[12:2] ? 10'h2ee : _GEN_1587; // @[Multiplier.scala 64:55]
  assign _GEN_1589 = 11'h635 == fractionSum[12:2] ? 10'h2ef : _GEN_1588; // @[Multiplier.scala 64:55]
  assign _GEN_1590 = 11'h636 == fractionSum[12:2] ? 10'h2ef : _GEN_1589; // @[Multiplier.scala 64:55]
  assign _GEN_1591 = 11'h637 == fractionSum[12:2] ? 10'h2f0 : _GEN_1590; // @[Multiplier.scala 64:55]
  assign _GEN_1592 = 11'h638 == fractionSum[12:2] ? 10'h2f0 : _GEN_1591; // @[Multiplier.scala 64:55]
  assign _GEN_1593 = 11'h639 == fractionSum[12:2] ? 10'h2f1 : _GEN_1592; // @[Multiplier.scala 64:55]
  assign _GEN_1594 = 11'h63a == fractionSum[12:2] ? 10'h2f1 : _GEN_1593; // @[Multiplier.scala 64:55]
  assign _GEN_1595 = 11'h63b == fractionSum[12:2] ? 10'h2f2 : _GEN_1594; // @[Multiplier.scala 64:55]
  assign _GEN_1596 = 11'h63c == fractionSum[12:2] ? 10'h2f2 : _GEN_1595; // @[Multiplier.scala 64:55]
  assign _GEN_1597 = 11'h63d == fractionSum[12:2] ? 10'h2f3 : _GEN_1596; // @[Multiplier.scala 64:55]
  assign _GEN_1598 = 11'h63e == fractionSum[12:2] ? 10'h2f3 : _GEN_1597; // @[Multiplier.scala 64:55]
  assign _GEN_1599 = 11'h63f == fractionSum[12:2] ? 10'h2f4 : _GEN_1598; // @[Multiplier.scala 64:55]
  assign _GEN_1600 = 11'h640 == fractionSum[12:2] ? 10'h2f4 : _GEN_1599; // @[Multiplier.scala 64:55]
  assign _GEN_1601 = 11'h641 == fractionSum[12:2] ? 10'h2f5 : _GEN_1600; // @[Multiplier.scala 64:55]
  assign _GEN_1602 = 11'h642 == fractionSum[12:2] ? 10'h2f5 : _GEN_1601; // @[Multiplier.scala 64:55]
  assign _GEN_1603 = 11'h643 == fractionSum[12:2] ? 10'h2f6 : _GEN_1602; // @[Multiplier.scala 64:55]
  assign _GEN_1604 = 11'h644 == fractionSum[12:2] ? 10'h2f6 : _GEN_1603; // @[Multiplier.scala 64:55]
  assign _GEN_1605 = 11'h645 == fractionSum[12:2] ? 10'h2f7 : _GEN_1604; // @[Multiplier.scala 64:55]
  assign _GEN_1606 = 11'h646 == fractionSum[12:2] ? 10'h2f7 : _GEN_1605; // @[Multiplier.scala 64:55]
  assign _GEN_1607 = 11'h647 == fractionSum[12:2] ? 10'h2f8 : _GEN_1606; // @[Multiplier.scala 64:55]
  assign _GEN_1608 = 11'h648 == fractionSum[12:2] ? 10'h2f8 : _GEN_1607; // @[Multiplier.scala 64:55]
  assign _GEN_1609 = 11'h649 == fractionSum[12:2] ? 10'h2f9 : _GEN_1608; // @[Multiplier.scala 64:55]
  assign _GEN_1610 = 11'h64a == fractionSum[12:2] ? 10'h2f9 : _GEN_1609; // @[Multiplier.scala 64:55]
  assign _GEN_1611 = 11'h64b == fractionSum[12:2] ? 10'h2fa : _GEN_1610; // @[Multiplier.scala 64:55]
  assign _GEN_1612 = 11'h64c == fractionSum[12:2] ? 10'h2fa : _GEN_1611; // @[Multiplier.scala 64:55]
  assign _GEN_1613 = 11'h64d == fractionSum[12:2] ? 10'h2fb : _GEN_1612; // @[Multiplier.scala 64:55]
  assign _GEN_1614 = 11'h64e == fractionSum[12:2] ? 10'h2fb : _GEN_1613; // @[Multiplier.scala 64:55]
  assign _GEN_1615 = 11'h64f == fractionSum[12:2] ? 10'h2fc : _GEN_1614; // @[Multiplier.scala 64:55]
  assign _GEN_1616 = 11'h650 == fractionSum[12:2] ? 10'h2fc : _GEN_1615; // @[Multiplier.scala 64:55]
  assign _GEN_1617 = 11'h651 == fractionSum[12:2] ? 10'h2fd : _GEN_1616; // @[Multiplier.scala 64:55]
  assign _GEN_1618 = 11'h652 == fractionSum[12:2] ? 10'h2fd : _GEN_1617; // @[Multiplier.scala 64:55]
  assign _GEN_1619 = 11'h653 == fractionSum[12:2] ? 10'h2fe : _GEN_1618; // @[Multiplier.scala 64:55]
  assign _GEN_1620 = 11'h654 == fractionSum[12:2] ? 10'h2fe : _GEN_1619; // @[Multiplier.scala 64:55]
  assign _GEN_1621 = 11'h655 == fractionSum[12:2] ? 10'h2ff : _GEN_1620; // @[Multiplier.scala 64:55]
  assign _GEN_1622 = 11'h656 == fractionSum[12:2] ? 10'h2ff : _GEN_1621; // @[Multiplier.scala 64:55]
  assign _GEN_1623 = 11'h657 == fractionSum[12:2] ? 10'h300 : _GEN_1622; // @[Multiplier.scala 64:55]
  assign _GEN_1624 = 11'h658 == fractionSum[12:2] ? 10'h301 : _GEN_1623; // @[Multiplier.scala 64:55]
  assign _GEN_1625 = 11'h659 == fractionSum[12:2] ? 10'h301 : _GEN_1624; // @[Multiplier.scala 64:55]
  assign _GEN_1626 = 11'h65a == fractionSum[12:2] ? 10'h302 : _GEN_1625; // @[Multiplier.scala 64:55]
  assign _GEN_1627 = 11'h65b == fractionSum[12:2] ? 10'h302 : _GEN_1626; // @[Multiplier.scala 64:55]
  assign _GEN_1628 = 11'h65c == fractionSum[12:2] ? 10'h303 : _GEN_1627; // @[Multiplier.scala 64:55]
  assign _GEN_1629 = 11'h65d == fractionSum[12:2] ? 10'h303 : _GEN_1628; // @[Multiplier.scala 64:55]
  assign _GEN_1630 = 11'h65e == fractionSum[12:2] ? 10'h304 : _GEN_1629; // @[Multiplier.scala 64:55]
  assign _GEN_1631 = 11'h65f == fractionSum[12:2] ? 10'h304 : _GEN_1630; // @[Multiplier.scala 64:55]
  assign _GEN_1632 = 11'h660 == fractionSum[12:2] ? 10'h305 : _GEN_1631; // @[Multiplier.scala 64:55]
  assign _GEN_1633 = 11'h661 == fractionSum[12:2] ? 10'h305 : _GEN_1632; // @[Multiplier.scala 64:55]
  assign _GEN_1634 = 11'h662 == fractionSum[12:2] ? 10'h306 : _GEN_1633; // @[Multiplier.scala 64:55]
  assign _GEN_1635 = 11'h663 == fractionSum[12:2] ? 10'h306 : _GEN_1634; // @[Multiplier.scala 64:55]
  assign _GEN_1636 = 11'h664 == fractionSum[12:2] ? 10'h307 : _GEN_1635; // @[Multiplier.scala 64:55]
  assign _GEN_1637 = 11'h665 == fractionSum[12:2] ? 10'h307 : _GEN_1636; // @[Multiplier.scala 64:55]
  assign _GEN_1638 = 11'h666 == fractionSum[12:2] ? 10'h308 : _GEN_1637; // @[Multiplier.scala 64:55]
  assign _GEN_1639 = 11'h667 == fractionSum[12:2] ? 10'h308 : _GEN_1638; // @[Multiplier.scala 64:55]
  assign _GEN_1640 = 11'h668 == fractionSum[12:2] ? 10'h309 : _GEN_1639; // @[Multiplier.scala 64:55]
  assign _GEN_1641 = 11'h669 == fractionSum[12:2] ? 10'h309 : _GEN_1640; // @[Multiplier.scala 64:55]
  assign _GEN_1642 = 11'h66a == fractionSum[12:2] ? 10'h30a : _GEN_1641; // @[Multiplier.scala 64:55]
  assign _GEN_1643 = 11'h66b == fractionSum[12:2] ? 10'h30a : _GEN_1642; // @[Multiplier.scala 64:55]
  assign _GEN_1644 = 11'h66c == fractionSum[12:2] ? 10'h30b : _GEN_1643; // @[Multiplier.scala 64:55]
  assign _GEN_1645 = 11'h66d == fractionSum[12:2] ? 10'h30c : _GEN_1644; // @[Multiplier.scala 64:55]
  assign _GEN_1646 = 11'h66e == fractionSum[12:2] ? 10'h30c : _GEN_1645; // @[Multiplier.scala 64:55]
  assign _GEN_1647 = 11'h66f == fractionSum[12:2] ? 10'h30d : _GEN_1646; // @[Multiplier.scala 64:55]
  assign _GEN_1648 = 11'h670 == fractionSum[12:2] ? 10'h30d : _GEN_1647; // @[Multiplier.scala 64:55]
  assign _GEN_1649 = 11'h671 == fractionSum[12:2] ? 10'h30e : _GEN_1648; // @[Multiplier.scala 64:55]
  assign _GEN_1650 = 11'h672 == fractionSum[12:2] ? 10'h30e : _GEN_1649; // @[Multiplier.scala 64:55]
  assign _GEN_1651 = 11'h673 == fractionSum[12:2] ? 10'h30f : _GEN_1650; // @[Multiplier.scala 64:55]
  assign _GEN_1652 = 11'h674 == fractionSum[12:2] ? 10'h30f : _GEN_1651; // @[Multiplier.scala 64:55]
  assign _GEN_1653 = 11'h675 == fractionSum[12:2] ? 10'h310 : _GEN_1652; // @[Multiplier.scala 64:55]
  assign _GEN_1654 = 11'h676 == fractionSum[12:2] ? 10'h310 : _GEN_1653; // @[Multiplier.scala 64:55]
  assign _GEN_1655 = 11'h677 == fractionSum[12:2] ? 10'h311 : _GEN_1654; // @[Multiplier.scala 64:55]
  assign _GEN_1656 = 11'h678 == fractionSum[12:2] ? 10'h311 : _GEN_1655; // @[Multiplier.scala 64:55]
  assign _GEN_1657 = 11'h679 == fractionSum[12:2] ? 10'h312 : _GEN_1656; // @[Multiplier.scala 64:55]
  assign _GEN_1658 = 11'h67a == fractionSum[12:2] ? 10'h312 : _GEN_1657; // @[Multiplier.scala 64:55]
  assign _GEN_1659 = 11'h67b == fractionSum[12:2] ? 10'h313 : _GEN_1658; // @[Multiplier.scala 64:55]
  assign _GEN_1660 = 11'h67c == fractionSum[12:2] ? 10'h313 : _GEN_1659; // @[Multiplier.scala 64:55]
  assign _GEN_1661 = 11'h67d == fractionSum[12:2] ? 10'h314 : _GEN_1660; // @[Multiplier.scala 64:55]
  assign _GEN_1662 = 11'h67e == fractionSum[12:2] ? 10'h315 : _GEN_1661; // @[Multiplier.scala 64:55]
  assign _GEN_1663 = 11'h67f == fractionSum[12:2] ? 10'h315 : _GEN_1662; // @[Multiplier.scala 64:55]
  assign _GEN_1664 = 11'h680 == fractionSum[12:2] ? 10'h316 : _GEN_1663; // @[Multiplier.scala 64:55]
  assign _GEN_1665 = 11'h681 == fractionSum[12:2] ? 10'h316 : _GEN_1664; // @[Multiplier.scala 64:55]
  assign _GEN_1666 = 11'h682 == fractionSum[12:2] ? 10'h317 : _GEN_1665; // @[Multiplier.scala 64:55]
  assign _GEN_1667 = 11'h683 == fractionSum[12:2] ? 10'h317 : _GEN_1666; // @[Multiplier.scala 64:55]
  assign _GEN_1668 = 11'h684 == fractionSum[12:2] ? 10'h318 : _GEN_1667; // @[Multiplier.scala 64:55]
  assign _GEN_1669 = 11'h685 == fractionSum[12:2] ? 10'h318 : _GEN_1668; // @[Multiplier.scala 64:55]
  assign _GEN_1670 = 11'h686 == fractionSum[12:2] ? 10'h319 : _GEN_1669; // @[Multiplier.scala 64:55]
  assign _GEN_1671 = 11'h687 == fractionSum[12:2] ? 10'h319 : _GEN_1670; // @[Multiplier.scala 64:55]
  assign _GEN_1672 = 11'h688 == fractionSum[12:2] ? 10'h31a : _GEN_1671; // @[Multiplier.scala 64:55]
  assign _GEN_1673 = 11'h689 == fractionSum[12:2] ? 10'h31a : _GEN_1672; // @[Multiplier.scala 64:55]
  assign _GEN_1674 = 11'h68a == fractionSum[12:2] ? 10'h31b : _GEN_1673; // @[Multiplier.scala 64:55]
  assign _GEN_1675 = 11'h68b == fractionSum[12:2] ? 10'h31c : _GEN_1674; // @[Multiplier.scala 64:55]
  assign _GEN_1676 = 11'h68c == fractionSum[12:2] ? 10'h31c : _GEN_1675; // @[Multiplier.scala 64:55]
  assign _GEN_1677 = 11'h68d == fractionSum[12:2] ? 10'h31d : _GEN_1676; // @[Multiplier.scala 64:55]
  assign _GEN_1678 = 11'h68e == fractionSum[12:2] ? 10'h31d : _GEN_1677; // @[Multiplier.scala 64:55]
  assign _GEN_1679 = 11'h68f == fractionSum[12:2] ? 10'h31e : _GEN_1678; // @[Multiplier.scala 64:55]
  assign _GEN_1680 = 11'h690 == fractionSum[12:2] ? 10'h31e : _GEN_1679; // @[Multiplier.scala 64:55]
  assign _GEN_1681 = 11'h691 == fractionSum[12:2] ? 10'h31f : _GEN_1680; // @[Multiplier.scala 64:55]
  assign _GEN_1682 = 11'h692 == fractionSum[12:2] ? 10'h31f : _GEN_1681; // @[Multiplier.scala 64:55]
  assign _GEN_1683 = 11'h693 == fractionSum[12:2] ? 10'h320 : _GEN_1682; // @[Multiplier.scala 64:55]
  assign _GEN_1684 = 11'h694 == fractionSum[12:2] ? 10'h320 : _GEN_1683; // @[Multiplier.scala 64:55]
  assign _GEN_1685 = 11'h695 == fractionSum[12:2] ? 10'h321 : _GEN_1684; // @[Multiplier.scala 64:55]
  assign _GEN_1686 = 11'h696 == fractionSum[12:2] ? 10'h321 : _GEN_1685; // @[Multiplier.scala 64:55]
  assign _GEN_1687 = 11'h697 == fractionSum[12:2] ? 10'h322 : _GEN_1686; // @[Multiplier.scala 64:55]
  assign _GEN_1688 = 11'h698 == fractionSum[12:2] ? 10'h323 : _GEN_1687; // @[Multiplier.scala 64:55]
  assign _GEN_1689 = 11'h699 == fractionSum[12:2] ? 10'h323 : _GEN_1688; // @[Multiplier.scala 64:55]
  assign _GEN_1690 = 11'h69a == fractionSum[12:2] ? 10'h324 : _GEN_1689; // @[Multiplier.scala 64:55]
  assign _GEN_1691 = 11'h69b == fractionSum[12:2] ? 10'h324 : _GEN_1690; // @[Multiplier.scala 64:55]
  assign _GEN_1692 = 11'h69c == fractionSum[12:2] ? 10'h325 : _GEN_1691; // @[Multiplier.scala 64:55]
  assign _GEN_1693 = 11'h69d == fractionSum[12:2] ? 10'h325 : _GEN_1692; // @[Multiplier.scala 64:55]
  assign _GEN_1694 = 11'h69e == fractionSum[12:2] ? 10'h326 : _GEN_1693; // @[Multiplier.scala 64:55]
  assign _GEN_1695 = 11'h69f == fractionSum[12:2] ? 10'h326 : _GEN_1694; // @[Multiplier.scala 64:55]
  assign _GEN_1696 = 11'h6a0 == fractionSum[12:2] ? 10'h327 : _GEN_1695; // @[Multiplier.scala 64:55]
  assign _GEN_1697 = 11'h6a1 == fractionSum[12:2] ? 10'h327 : _GEN_1696; // @[Multiplier.scala 64:55]
  assign _GEN_1698 = 11'h6a2 == fractionSum[12:2] ? 10'h328 : _GEN_1697; // @[Multiplier.scala 64:55]
  assign _GEN_1699 = 11'h6a3 == fractionSum[12:2] ? 10'h329 : _GEN_1698; // @[Multiplier.scala 64:55]
  assign _GEN_1700 = 11'h6a4 == fractionSum[12:2] ? 10'h329 : _GEN_1699; // @[Multiplier.scala 64:55]
  assign _GEN_1701 = 11'h6a5 == fractionSum[12:2] ? 10'h32a : _GEN_1700; // @[Multiplier.scala 64:55]
  assign _GEN_1702 = 11'h6a6 == fractionSum[12:2] ? 10'h32a : _GEN_1701; // @[Multiplier.scala 64:55]
  assign _GEN_1703 = 11'h6a7 == fractionSum[12:2] ? 10'h32b : _GEN_1702; // @[Multiplier.scala 64:55]
  assign _GEN_1704 = 11'h6a8 == fractionSum[12:2] ? 10'h32b : _GEN_1703; // @[Multiplier.scala 64:55]
  assign _GEN_1705 = 11'h6a9 == fractionSum[12:2] ? 10'h32c : _GEN_1704; // @[Multiplier.scala 64:55]
  assign _GEN_1706 = 11'h6aa == fractionSum[12:2] ? 10'h32c : _GEN_1705; // @[Multiplier.scala 64:55]
  assign _GEN_1707 = 11'h6ab == fractionSum[12:2] ? 10'h32d : _GEN_1706; // @[Multiplier.scala 64:55]
  assign _GEN_1708 = 11'h6ac == fractionSum[12:2] ? 10'h32d : _GEN_1707; // @[Multiplier.scala 64:55]
  assign _GEN_1709 = 11'h6ad == fractionSum[12:2] ? 10'h32e : _GEN_1708; // @[Multiplier.scala 64:55]
  assign _GEN_1710 = 11'h6ae == fractionSum[12:2] ? 10'h32f : _GEN_1709; // @[Multiplier.scala 64:55]
  assign _GEN_1711 = 11'h6af == fractionSum[12:2] ? 10'h32f : _GEN_1710; // @[Multiplier.scala 64:55]
  assign _GEN_1712 = 11'h6b0 == fractionSum[12:2] ? 10'h330 : _GEN_1711; // @[Multiplier.scala 64:55]
  assign _GEN_1713 = 11'h6b1 == fractionSum[12:2] ? 10'h330 : _GEN_1712; // @[Multiplier.scala 64:55]
  assign _GEN_1714 = 11'h6b2 == fractionSum[12:2] ? 10'h331 : _GEN_1713; // @[Multiplier.scala 64:55]
  assign _GEN_1715 = 11'h6b3 == fractionSum[12:2] ? 10'h331 : _GEN_1714; // @[Multiplier.scala 64:55]
  assign _GEN_1716 = 11'h6b4 == fractionSum[12:2] ? 10'h332 : _GEN_1715; // @[Multiplier.scala 64:55]
  assign _GEN_1717 = 11'h6b5 == fractionSum[12:2] ? 10'h332 : _GEN_1716; // @[Multiplier.scala 64:55]
  assign _GEN_1718 = 11'h6b6 == fractionSum[12:2] ? 10'h333 : _GEN_1717; // @[Multiplier.scala 64:55]
  assign _GEN_1719 = 11'h6b7 == fractionSum[12:2] ? 10'h334 : _GEN_1718; // @[Multiplier.scala 64:55]
  assign _GEN_1720 = 11'h6b8 == fractionSum[12:2] ? 10'h334 : _GEN_1719; // @[Multiplier.scala 64:55]
  assign _GEN_1721 = 11'h6b9 == fractionSum[12:2] ? 10'h335 : _GEN_1720; // @[Multiplier.scala 64:55]
  assign _GEN_1722 = 11'h6ba == fractionSum[12:2] ? 10'h335 : _GEN_1721; // @[Multiplier.scala 64:55]
  assign _GEN_1723 = 11'h6bb == fractionSum[12:2] ? 10'h336 : _GEN_1722; // @[Multiplier.scala 64:55]
  assign _GEN_1724 = 11'h6bc == fractionSum[12:2] ? 10'h336 : _GEN_1723; // @[Multiplier.scala 64:55]
  assign _GEN_1725 = 11'h6bd == fractionSum[12:2] ? 10'h337 : _GEN_1724; // @[Multiplier.scala 64:55]
  assign _GEN_1726 = 11'h6be == fractionSum[12:2] ? 10'h337 : _GEN_1725; // @[Multiplier.scala 64:55]
  assign _GEN_1727 = 11'h6bf == fractionSum[12:2] ? 10'h338 : _GEN_1726; // @[Multiplier.scala 64:55]
  assign _GEN_1728 = 11'h6c0 == fractionSum[12:2] ? 10'h339 : _GEN_1727; // @[Multiplier.scala 64:55]
  assign _GEN_1729 = 11'h6c1 == fractionSum[12:2] ? 10'h339 : _GEN_1728; // @[Multiplier.scala 64:55]
  assign _GEN_1730 = 11'h6c2 == fractionSum[12:2] ? 10'h33a : _GEN_1729; // @[Multiplier.scala 64:55]
  assign _GEN_1731 = 11'h6c3 == fractionSum[12:2] ? 10'h33a : _GEN_1730; // @[Multiplier.scala 64:55]
  assign _GEN_1732 = 11'h6c4 == fractionSum[12:2] ? 10'h33b : _GEN_1731; // @[Multiplier.scala 64:55]
  assign _GEN_1733 = 11'h6c5 == fractionSum[12:2] ? 10'h33b : _GEN_1732; // @[Multiplier.scala 64:55]
  assign _GEN_1734 = 11'h6c6 == fractionSum[12:2] ? 10'h33c : _GEN_1733; // @[Multiplier.scala 64:55]
  assign _GEN_1735 = 11'h6c7 == fractionSum[12:2] ? 10'h33c : _GEN_1734; // @[Multiplier.scala 64:55]
  assign _GEN_1736 = 11'h6c8 == fractionSum[12:2] ? 10'h33d : _GEN_1735; // @[Multiplier.scala 64:55]
  assign _GEN_1737 = 11'h6c9 == fractionSum[12:2] ? 10'h33e : _GEN_1736; // @[Multiplier.scala 64:55]
  assign _GEN_1738 = 11'h6ca == fractionSum[12:2] ? 10'h33e : _GEN_1737; // @[Multiplier.scala 64:55]
  assign _GEN_1739 = 11'h6cb == fractionSum[12:2] ? 10'h33f : _GEN_1738; // @[Multiplier.scala 64:55]
  assign _GEN_1740 = 11'h6cc == fractionSum[12:2] ? 10'h33f : _GEN_1739; // @[Multiplier.scala 64:55]
  assign _GEN_1741 = 11'h6cd == fractionSum[12:2] ? 10'h340 : _GEN_1740; // @[Multiplier.scala 64:55]
  assign _GEN_1742 = 11'h6ce == fractionSum[12:2] ? 10'h340 : _GEN_1741; // @[Multiplier.scala 64:55]
  assign _GEN_1743 = 11'h6cf == fractionSum[12:2] ? 10'h341 : _GEN_1742; // @[Multiplier.scala 64:55]
  assign _GEN_1744 = 11'h6d0 == fractionSum[12:2] ? 10'h342 : _GEN_1743; // @[Multiplier.scala 64:55]
  assign _GEN_1745 = 11'h6d1 == fractionSum[12:2] ? 10'h342 : _GEN_1744; // @[Multiplier.scala 64:55]
  assign _GEN_1746 = 11'h6d2 == fractionSum[12:2] ? 10'h343 : _GEN_1745; // @[Multiplier.scala 64:55]
  assign _GEN_1747 = 11'h6d3 == fractionSum[12:2] ? 10'h343 : _GEN_1746; // @[Multiplier.scala 64:55]
  assign _GEN_1748 = 11'h6d4 == fractionSum[12:2] ? 10'h344 : _GEN_1747; // @[Multiplier.scala 64:55]
  assign _GEN_1749 = 11'h6d5 == fractionSum[12:2] ? 10'h344 : _GEN_1748; // @[Multiplier.scala 64:55]
  assign _GEN_1750 = 11'h6d6 == fractionSum[12:2] ? 10'h345 : _GEN_1749; // @[Multiplier.scala 64:55]
  assign _GEN_1751 = 11'h6d7 == fractionSum[12:2] ? 10'h346 : _GEN_1750; // @[Multiplier.scala 64:55]
  assign _GEN_1752 = 11'h6d8 == fractionSum[12:2] ? 10'h346 : _GEN_1751; // @[Multiplier.scala 64:55]
  assign _GEN_1753 = 11'h6d9 == fractionSum[12:2] ? 10'h347 : _GEN_1752; // @[Multiplier.scala 64:55]
  assign _GEN_1754 = 11'h6da == fractionSum[12:2] ? 10'h347 : _GEN_1753; // @[Multiplier.scala 64:55]
  assign _GEN_1755 = 11'h6db == fractionSum[12:2] ? 10'h348 : _GEN_1754; // @[Multiplier.scala 64:55]
  assign _GEN_1756 = 11'h6dc == fractionSum[12:2] ? 10'h348 : _GEN_1755; // @[Multiplier.scala 64:55]
  assign _GEN_1757 = 11'h6dd == fractionSum[12:2] ? 10'h349 : _GEN_1756; // @[Multiplier.scala 64:55]
  assign _GEN_1758 = 11'h6de == fractionSum[12:2] ? 10'h349 : _GEN_1757; // @[Multiplier.scala 64:55]
  assign _GEN_1759 = 11'h6df == fractionSum[12:2] ? 10'h34a : _GEN_1758; // @[Multiplier.scala 64:55]
  assign _GEN_1760 = 11'h6e0 == fractionSum[12:2] ? 10'h34b : _GEN_1759; // @[Multiplier.scala 64:55]
  assign _GEN_1761 = 11'h6e1 == fractionSum[12:2] ? 10'h34b : _GEN_1760; // @[Multiplier.scala 64:55]
  assign _GEN_1762 = 11'h6e2 == fractionSum[12:2] ? 10'h34c : _GEN_1761; // @[Multiplier.scala 64:55]
  assign _GEN_1763 = 11'h6e3 == fractionSum[12:2] ? 10'h34c : _GEN_1762; // @[Multiplier.scala 64:55]
  assign _GEN_1764 = 11'h6e4 == fractionSum[12:2] ? 10'h34d : _GEN_1763; // @[Multiplier.scala 64:55]
  assign _GEN_1765 = 11'h6e5 == fractionSum[12:2] ? 10'h34d : _GEN_1764; // @[Multiplier.scala 64:55]
  assign _GEN_1766 = 11'h6e6 == fractionSum[12:2] ? 10'h34e : _GEN_1765; // @[Multiplier.scala 64:55]
  assign _GEN_1767 = 11'h6e7 == fractionSum[12:2] ? 10'h34f : _GEN_1766; // @[Multiplier.scala 64:55]
  assign _GEN_1768 = 11'h6e8 == fractionSum[12:2] ? 10'h34f : _GEN_1767; // @[Multiplier.scala 64:55]
  assign _GEN_1769 = 11'h6e9 == fractionSum[12:2] ? 10'h350 : _GEN_1768; // @[Multiplier.scala 64:55]
  assign _GEN_1770 = 11'h6ea == fractionSum[12:2] ? 10'h350 : _GEN_1769; // @[Multiplier.scala 64:55]
  assign _GEN_1771 = 11'h6eb == fractionSum[12:2] ? 10'h351 : _GEN_1770; // @[Multiplier.scala 64:55]
  assign _GEN_1772 = 11'h6ec == fractionSum[12:2] ? 10'h351 : _GEN_1771; // @[Multiplier.scala 64:55]
  assign _GEN_1773 = 11'h6ed == fractionSum[12:2] ? 10'h352 : _GEN_1772; // @[Multiplier.scala 64:55]
  assign _GEN_1774 = 11'h6ee == fractionSum[12:2] ? 10'h353 : _GEN_1773; // @[Multiplier.scala 64:55]
  assign _GEN_1775 = 11'h6ef == fractionSum[12:2] ? 10'h353 : _GEN_1774; // @[Multiplier.scala 64:55]
  assign _GEN_1776 = 11'h6f0 == fractionSum[12:2] ? 10'h354 : _GEN_1775; // @[Multiplier.scala 64:55]
  assign _GEN_1777 = 11'h6f1 == fractionSum[12:2] ? 10'h354 : _GEN_1776; // @[Multiplier.scala 64:55]
  assign _GEN_1778 = 11'h6f2 == fractionSum[12:2] ? 10'h355 : _GEN_1777; // @[Multiplier.scala 64:55]
  assign _GEN_1779 = 11'h6f3 == fractionSum[12:2] ? 10'h356 : _GEN_1778; // @[Multiplier.scala 64:55]
  assign _GEN_1780 = 11'h6f4 == fractionSum[12:2] ? 10'h356 : _GEN_1779; // @[Multiplier.scala 64:55]
  assign _GEN_1781 = 11'h6f5 == fractionSum[12:2] ? 10'h357 : _GEN_1780; // @[Multiplier.scala 64:55]
  assign _GEN_1782 = 11'h6f6 == fractionSum[12:2] ? 10'h357 : _GEN_1781; // @[Multiplier.scala 64:55]
  assign _GEN_1783 = 11'h6f7 == fractionSum[12:2] ? 10'h358 : _GEN_1782; // @[Multiplier.scala 64:55]
  assign _GEN_1784 = 11'h6f8 == fractionSum[12:2] ? 10'h358 : _GEN_1783; // @[Multiplier.scala 64:55]
  assign _GEN_1785 = 11'h6f9 == fractionSum[12:2] ? 10'h359 : _GEN_1784; // @[Multiplier.scala 64:55]
  assign _GEN_1786 = 11'h6fa == fractionSum[12:2] ? 10'h35a : _GEN_1785; // @[Multiplier.scala 64:55]
  assign _GEN_1787 = 11'h6fb == fractionSum[12:2] ? 10'h35a : _GEN_1786; // @[Multiplier.scala 64:55]
  assign _GEN_1788 = 11'h6fc == fractionSum[12:2] ? 10'h35b : _GEN_1787; // @[Multiplier.scala 64:55]
  assign _GEN_1789 = 11'h6fd == fractionSum[12:2] ? 10'h35b : _GEN_1788; // @[Multiplier.scala 64:55]
  assign _GEN_1790 = 11'h6fe == fractionSum[12:2] ? 10'h35c : _GEN_1789; // @[Multiplier.scala 64:55]
  assign _GEN_1791 = 11'h6ff == fractionSum[12:2] ? 10'h35c : _GEN_1790; // @[Multiplier.scala 64:55]
  assign _GEN_1792 = 11'h700 == fractionSum[12:2] ? 10'h35d : _GEN_1791; // @[Multiplier.scala 64:55]
  assign _GEN_1793 = 11'h701 == fractionSum[12:2] ? 10'h35e : _GEN_1792; // @[Multiplier.scala 64:55]
  assign _GEN_1794 = 11'h702 == fractionSum[12:2] ? 10'h35e : _GEN_1793; // @[Multiplier.scala 64:55]
  assign _GEN_1795 = 11'h703 == fractionSum[12:2] ? 10'h35f : _GEN_1794; // @[Multiplier.scala 64:55]
  assign _GEN_1796 = 11'h704 == fractionSum[12:2] ? 10'h35f : _GEN_1795; // @[Multiplier.scala 64:55]
  assign _GEN_1797 = 11'h705 == fractionSum[12:2] ? 10'h360 : _GEN_1796; // @[Multiplier.scala 64:55]
  assign _GEN_1798 = 11'h706 == fractionSum[12:2] ? 10'h361 : _GEN_1797; // @[Multiplier.scala 64:55]
  assign _GEN_1799 = 11'h707 == fractionSum[12:2] ? 10'h361 : _GEN_1798; // @[Multiplier.scala 64:55]
  assign _GEN_1800 = 11'h708 == fractionSum[12:2] ? 10'h362 : _GEN_1799; // @[Multiplier.scala 64:55]
  assign _GEN_1801 = 11'h709 == fractionSum[12:2] ? 10'h362 : _GEN_1800; // @[Multiplier.scala 64:55]
  assign _GEN_1802 = 11'h70a == fractionSum[12:2] ? 10'h363 : _GEN_1801; // @[Multiplier.scala 64:55]
  assign _GEN_1803 = 11'h70b == fractionSum[12:2] ? 10'h364 : _GEN_1802; // @[Multiplier.scala 64:55]
  assign _GEN_1804 = 11'h70c == fractionSum[12:2] ? 10'h364 : _GEN_1803; // @[Multiplier.scala 64:55]
  assign _GEN_1805 = 11'h70d == fractionSum[12:2] ? 10'h365 : _GEN_1804; // @[Multiplier.scala 64:55]
  assign _GEN_1806 = 11'h70e == fractionSum[12:2] ? 10'h365 : _GEN_1805; // @[Multiplier.scala 64:55]
  assign _GEN_1807 = 11'h70f == fractionSum[12:2] ? 10'h366 : _GEN_1806; // @[Multiplier.scala 64:55]
  assign _GEN_1808 = 11'h710 == fractionSum[12:2] ? 10'h366 : _GEN_1807; // @[Multiplier.scala 64:55]
  assign _GEN_1809 = 11'h711 == fractionSum[12:2] ? 10'h367 : _GEN_1808; // @[Multiplier.scala 64:55]
  assign _GEN_1810 = 11'h712 == fractionSum[12:2] ? 10'h368 : _GEN_1809; // @[Multiplier.scala 64:55]
  assign _GEN_1811 = 11'h713 == fractionSum[12:2] ? 10'h368 : _GEN_1810; // @[Multiplier.scala 64:55]
  assign _GEN_1812 = 11'h714 == fractionSum[12:2] ? 10'h369 : _GEN_1811; // @[Multiplier.scala 64:55]
  assign _GEN_1813 = 11'h715 == fractionSum[12:2] ? 10'h369 : _GEN_1812; // @[Multiplier.scala 64:55]
  assign _GEN_1814 = 11'h716 == fractionSum[12:2] ? 10'h36a : _GEN_1813; // @[Multiplier.scala 64:55]
  assign _GEN_1815 = 11'h717 == fractionSum[12:2] ? 10'h36b : _GEN_1814; // @[Multiplier.scala 64:55]
  assign _GEN_1816 = 11'h718 == fractionSum[12:2] ? 10'h36b : _GEN_1815; // @[Multiplier.scala 64:55]
  assign _GEN_1817 = 11'h719 == fractionSum[12:2] ? 10'h36c : _GEN_1816; // @[Multiplier.scala 64:55]
  assign _GEN_1818 = 11'h71a == fractionSum[12:2] ? 10'h36c : _GEN_1817; // @[Multiplier.scala 64:55]
  assign _GEN_1819 = 11'h71b == fractionSum[12:2] ? 10'h36d : _GEN_1818; // @[Multiplier.scala 64:55]
  assign _GEN_1820 = 11'h71c == fractionSum[12:2] ? 10'h36e : _GEN_1819; // @[Multiplier.scala 64:55]
  assign _GEN_1821 = 11'h71d == fractionSum[12:2] ? 10'h36e : _GEN_1820; // @[Multiplier.scala 64:55]
  assign _GEN_1822 = 11'h71e == fractionSum[12:2] ? 10'h36f : _GEN_1821; // @[Multiplier.scala 64:55]
  assign _GEN_1823 = 11'h71f == fractionSum[12:2] ? 10'h36f : _GEN_1822; // @[Multiplier.scala 64:55]
  assign _GEN_1824 = 11'h720 == fractionSum[12:2] ? 10'h370 : _GEN_1823; // @[Multiplier.scala 64:55]
  assign _GEN_1825 = 11'h721 == fractionSum[12:2] ? 10'h371 : _GEN_1824; // @[Multiplier.scala 64:55]
  assign _GEN_1826 = 11'h722 == fractionSum[12:2] ? 10'h371 : _GEN_1825; // @[Multiplier.scala 64:55]
  assign _GEN_1827 = 11'h723 == fractionSum[12:2] ? 10'h372 : _GEN_1826; // @[Multiplier.scala 64:55]
  assign _GEN_1828 = 11'h724 == fractionSum[12:2] ? 10'h372 : _GEN_1827; // @[Multiplier.scala 64:55]
  assign _GEN_1829 = 11'h725 == fractionSum[12:2] ? 10'h373 : _GEN_1828; // @[Multiplier.scala 64:55]
  assign _GEN_1830 = 11'h726 == fractionSum[12:2] ? 10'h374 : _GEN_1829; // @[Multiplier.scala 64:55]
  assign _GEN_1831 = 11'h727 == fractionSum[12:2] ? 10'h374 : _GEN_1830; // @[Multiplier.scala 64:55]
  assign _GEN_1832 = 11'h728 == fractionSum[12:2] ? 10'h375 : _GEN_1831; // @[Multiplier.scala 64:55]
  assign _GEN_1833 = 11'h729 == fractionSum[12:2] ? 10'h375 : _GEN_1832; // @[Multiplier.scala 64:55]
  assign _GEN_1834 = 11'h72a == fractionSum[12:2] ? 10'h376 : _GEN_1833; // @[Multiplier.scala 64:55]
  assign _GEN_1835 = 11'h72b == fractionSum[12:2] ? 10'h377 : _GEN_1834; // @[Multiplier.scala 64:55]
  assign _GEN_1836 = 11'h72c == fractionSum[12:2] ? 10'h377 : _GEN_1835; // @[Multiplier.scala 64:55]
  assign _GEN_1837 = 11'h72d == fractionSum[12:2] ? 10'h378 : _GEN_1836; // @[Multiplier.scala 64:55]
  assign _GEN_1838 = 11'h72e == fractionSum[12:2] ? 10'h378 : _GEN_1837; // @[Multiplier.scala 64:55]
  assign _GEN_1839 = 11'h72f == fractionSum[12:2] ? 10'h379 : _GEN_1838; // @[Multiplier.scala 64:55]
  assign _GEN_1840 = 11'h730 == fractionSum[12:2] ? 10'h37a : _GEN_1839; // @[Multiplier.scala 64:55]
  assign _GEN_1841 = 11'h731 == fractionSum[12:2] ? 10'h37a : _GEN_1840; // @[Multiplier.scala 64:55]
  assign _GEN_1842 = 11'h732 == fractionSum[12:2] ? 10'h37b : _GEN_1841; // @[Multiplier.scala 64:55]
  assign _GEN_1843 = 11'h733 == fractionSum[12:2] ? 10'h37b : _GEN_1842; // @[Multiplier.scala 64:55]
  assign _GEN_1844 = 11'h734 == fractionSum[12:2] ? 10'h37c : _GEN_1843; // @[Multiplier.scala 64:55]
  assign _GEN_1845 = 11'h735 == fractionSum[12:2] ? 10'h37d : _GEN_1844; // @[Multiplier.scala 64:55]
  assign _GEN_1846 = 11'h736 == fractionSum[12:2] ? 10'h37d : _GEN_1845; // @[Multiplier.scala 64:55]
  assign _GEN_1847 = 11'h737 == fractionSum[12:2] ? 10'h37e : _GEN_1846; // @[Multiplier.scala 64:55]
  assign _GEN_1848 = 11'h738 == fractionSum[12:2] ? 10'h37e : _GEN_1847; // @[Multiplier.scala 64:55]
  assign _GEN_1849 = 11'h739 == fractionSum[12:2] ? 10'h37f : _GEN_1848; // @[Multiplier.scala 64:55]
  assign _GEN_1850 = 11'h73a == fractionSum[12:2] ? 10'h380 : _GEN_1849; // @[Multiplier.scala 64:55]
  assign _GEN_1851 = 11'h73b == fractionSum[12:2] ? 10'h380 : _GEN_1850; // @[Multiplier.scala 64:55]
  assign _GEN_1852 = 11'h73c == fractionSum[12:2] ? 10'h381 : _GEN_1851; // @[Multiplier.scala 64:55]
  assign _GEN_1853 = 11'h73d == fractionSum[12:2] ? 10'h381 : _GEN_1852; // @[Multiplier.scala 64:55]
  assign _GEN_1854 = 11'h73e == fractionSum[12:2] ? 10'h382 : _GEN_1853; // @[Multiplier.scala 64:55]
  assign _GEN_1855 = 11'h73f == fractionSum[12:2] ? 10'h383 : _GEN_1854; // @[Multiplier.scala 64:55]
  assign _GEN_1856 = 11'h740 == fractionSum[12:2] ? 10'h383 : _GEN_1855; // @[Multiplier.scala 64:55]
  assign _GEN_1857 = 11'h741 == fractionSum[12:2] ? 10'h384 : _GEN_1856; // @[Multiplier.scala 64:55]
  assign _GEN_1858 = 11'h742 == fractionSum[12:2] ? 10'h384 : _GEN_1857; // @[Multiplier.scala 64:55]
  assign _GEN_1859 = 11'h743 == fractionSum[12:2] ? 10'h385 : _GEN_1858; // @[Multiplier.scala 64:55]
  assign _GEN_1860 = 11'h744 == fractionSum[12:2] ? 10'h386 : _GEN_1859; // @[Multiplier.scala 64:55]
  assign _GEN_1861 = 11'h745 == fractionSum[12:2] ? 10'h386 : _GEN_1860; // @[Multiplier.scala 64:55]
  assign _GEN_1862 = 11'h746 == fractionSum[12:2] ? 10'h387 : _GEN_1861; // @[Multiplier.scala 64:55]
  assign _GEN_1863 = 11'h747 == fractionSum[12:2] ? 10'h387 : _GEN_1862; // @[Multiplier.scala 64:55]
  assign _GEN_1864 = 11'h748 == fractionSum[12:2] ? 10'h388 : _GEN_1863; // @[Multiplier.scala 64:55]
  assign _GEN_1865 = 11'h749 == fractionSum[12:2] ? 10'h389 : _GEN_1864; // @[Multiplier.scala 64:55]
  assign _GEN_1866 = 11'h74a == fractionSum[12:2] ? 10'h389 : _GEN_1865; // @[Multiplier.scala 64:55]
  assign _GEN_1867 = 11'h74b == fractionSum[12:2] ? 10'h38a : _GEN_1866; // @[Multiplier.scala 64:55]
  assign _GEN_1868 = 11'h74c == fractionSum[12:2] ? 10'h38b : _GEN_1867; // @[Multiplier.scala 64:55]
  assign _GEN_1869 = 11'h74d == fractionSum[12:2] ? 10'h38b : _GEN_1868; // @[Multiplier.scala 64:55]
  assign _GEN_1870 = 11'h74e == fractionSum[12:2] ? 10'h38c : _GEN_1869; // @[Multiplier.scala 64:55]
  assign _GEN_1871 = 11'h74f == fractionSum[12:2] ? 10'h38c : _GEN_1870; // @[Multiplier.scala 64:55]
  assign _GEN_1872 = 11'h750 == fractionSum[12:2] ? 10'h38d : _GEN_1871; // @[Multiplier.scala 64:55]
  assign _GEN_1873 = 11'h751 == fractionSum[12:2] ? 10'h38e : _GEN_1872; // @[Multiplier.scala 64:55]
  assign _GEN_1874 = 11'h752 == fractionSum[12:2] ? 10'h38e : _GEN_1873; // @[Multiplier.scala 64:55]
  assign _GEN_1875 = 11'h753 == fractionSum[12:2] ? 10'h38f : _GEN_1874; // @[Multiplier.scala 64:55]
  assign _GEN_1876 = 11'h754 == fractionSum[12:2] ? 10'h38f : _GEN_1875; // @[Multiplier.scala 64:55]
  assign _GEN_1877 = 11'h755 == fractionSum[12:2] ? 10'h390 : _GEN_1876; // @[Multiplier.scala 64:55]
  assign _GEN_1878 = 11'h756 == fractionSum[12:2] ? 10'h391 : _GEN_1877; // @[Multiplier.scala 64:55]
  assign _GEN_1879 = 11'h757 == fractionSum[12:2] ? 10'h391 : _GEN_1878; // @[Multiplier.scala 64:55]
  assign _GEN_1880 = 11'h758 == fractionSum[12:2] ? 10'h392 : _GEN_1879; // @[Multiplier.scala 64:55]
  assign _GEN_1881 = 11'h759 == fractionSum[12:2] ? 10'h393 : _GEN_1880; // @[Multiplier.scala 64:55]
  assign _GEN_1882 = 11'h75a == fractionSum[12:2] ? 10'h393 : _GEN_1881; // @[Multiplier.scala 64:55]
  assign _GEN_1883 = 11'h75b == fractionSum[12:2] ? 10'h394 : _GEN_1882; // @[Multiplier.scala 64:55]
  assign _GEN_1884 = 11'h75c == fractionSum[12:2] ? 10'h394 : _GEN_1883; // @[Multiplier.scala 64:55]
  assign _GEN_1885 = 11'h75d == fractionSum[12:2] ? 10'h395 : _GEN_1884; // @[Multiplier.scala 64:55]
  assign _GEN_1886 = 11'h75e == fractionSum[12:2] ? 10'h396 : _GEN_1885; // @[Multiplier.scala 64:55]
  assign _GEN_1887 = 11'h75f == fractionSum[12:2] ? 10'h396 : _GEN_1886; // @[Multiplier.scala 64:55]
  assign _GEN_1888 = 11'h760 == fractionSum[12:2] ? 10'h397 : _GEN_1887; // @[Multiplier.scala 64:55]
  assign _GEN_1889 = 11'h761 == fractionSum[12:2] ? 10'h398 : _GEN_1888; // @[Multiplier.scala 64:55]
  assign _GEN_1890 = 11'h762 == fractionSum[12:2] ? 10'h398 : _GEN_1889; // @[Multiplier.scala 64:55]
  assign _GEN_1891 = 11'h763 == fractionSum[12:2] ? 10'h399 : _GEN_1890; // @[Multiplier.scala 64:55]
  assign _GEN_1892 = 11'h764 == fractionSum[12:2] ? 10'h399 : _GEN_1891; // @[Multiplier.scala 64:55]
  assign _GEN_1893 = 11'h765 == fractionSum[12:2] ? 10'h39a : _GEN_1892; // @[Multiplier.scala 64:55]
  assign _GEN_1894 = 11'h766 == fractionSum[12:2] ? 10'h39b : _GEN_1893; // @[Multiplier.scala 64:55]
  assign _GEN_1895 = 11'h767 == fractionSum[12:2] ? 10'h39b : _GEN_1894; // @[Multiplier.scala 64:55]
  assign _GEN_1896 = 11'h768 == fractionSum[12:2] ? 10'h39c : _GEN_1895; // @[Multiplier.scala 64:55]
  assign _GEN_1897 = 11'h769 == fractionSum[12:2] ? 10'h39d : _GEN_1896; // @[Multiplier.scala 64:55]
  assign _GEN_1898 = 11'h76a == fractionSum[12:2] ? 10'h39d : _GEN_1897; // @[Multiplier.scala 64:55]
  assign _GEN_1899 = 11'h76b == fractionSum[12:2] ? 10'h39e : _GEN_1898; // @[Multiplier.scala 64:55]
  assign _GEN_1900 = 11'h76c == fractionSum[12:2] ? 10'h39e : _GEN_1899; // @[Multiplier.scala 64:55]
  assign _GEN_1901 = 11'h76d == fractionSum[12:2] ? 10'h39f : _GEN_1900; // @[Multiplier.scala 64:55]
  assign _GEN_1902 = 11'h76e == fractionSum[12:2] ? 10'h3a0 : _GEN_1901; // @[Multiplier.scala 64:55]
  assign _GEN_1903 = 11'h76f == fractionSum[12:2] ? 10'h3a0 : _GEN_1902; // @[Multiplier.scala 64:55]
  assign _GEN_1904 = 11'h770 == fractionSum[12:2] ? 10'h3a1 : _GEN_1903; // @[Multiplier.scala 64:55]
  assign _GEN_1905 = 11'h771 == fractionSum[12:2] ? 10'h3a2 : _GEN_1904; // @[Multiplier.scala 64:55]
  assign _GEN_1906 = 11'h772 == fractionSum[12:2] ? 10'h3a2 : _GEN_1905; // @[Multiplier.scala 64:55]
  assign _GEN_1907 = 11'h773 == fractionSum[12:2] ? 10'h3a3 : _GEN_1906; // @[Multiplier.scala 64:55]
  assign _GEN_1908 = 11'h774 == fractionSum[12:2] ? 10'h3a3 : _GEN_1907; // @[Multiplier.scala 64:55]
  assign _GEN_1909 = 11'h775 == fractionSum[12:2] ? 10'h3a4 : _GEN_1908; // @[Multiplier.scala 64:55]
  assign _GEN_1910 = 11'h776 == fractionSum[12:2] ? 10'h3a5 : _GEN_1909; // @[Multiplier.scala 64:55]
  assign _GEN_1911 = 11'h777 == fractionSum[12:2] ? 10'h3a5 : _GEN_1910; // @[Multiplier.scala 64:55]
  assign _GEN_1912 = 11'h778 == fractionSum[12:2] ? 10'h3a6 : _GEN_1911; // @[Multiplier.scala 64:55]
  assign _GEN_1913 = 11'h779 == fractionSum[12:2] ? 10'h3a7 : _GEN_1912; // @[Multiplier.scala 64:55]
  assign _GEN_1914 = 11'h77a == fractionSum[12:2] ? 10'h3a7 : _GEN_1913; // @[Multiplier.scala 64:55]
  assign _GEN_1915 = 11'h77b == fractionSum[12:2] ? 10'h3a8 : _GEN_1914; // @[Multiplier.scala 64:55]
  assign _GEN_1916 = 11'h77c == fractionSum[12:2] ? 10'h3a8 : _GEN_1915; // @[Multiplier.scala 64:55]
  assign _GEN_1917 = 11'h77d == fractionSum[12:2] ? 10'h3a9 : _GEN_1916; // @[Multiplier.scala 64:55]
  assign _GEN_1918 = 11'h77e == fractionSum[12:2] ? 10'h3aa : _GEN_1917; // @[Multiplier.scala 64:55]
  assign _GEN_1919 = 11'h77f == fractionSum[12:2] ? 10'h3aa : _GEN_1918; // @[Multiplier.scala 64:55]
  assign _GEN_1920 = 11'h780 == fractionSum[12:2] ? 10'h3ab : _GEN_1919; // @[Multiplier.scala 64:55]
  assign _GEN_1921 = 11'h781 == fractionSum[12:2] ? 10'h3ac : _GEN_1920; // @[Multiplier.scala 64:55]
  assign _GEN_1922 = 11'h782 == fractionSum[12:2] ? 10'h3ac : _GEN_1921; // @[Multiplier.scala 64:55]
  assign _GEN_1923 = 11'h783 == fractionSum[12:2] ? 10'h3ad : _GEN_1922; // @[Multiplier.scala 64:55]
  assign _GEN_1924 = 11'h784 == fractionSum[12:2] ? 10'h3ae : _GEN_1923; // @[Multiplier.scala 64:55]
  assign _GEN_1925 = 11'h785 == fractionSum[12:2] ? 10'h3ae : _GEN_1924; // @[Multiplier.scala 64:55]
  assign _GEN_1926 = 11'h786 == fractionSum[12:2] ? 10'h3af : _GEN_1925; // @[Multiplier.scala 64:55]
  assign _GEN_1927 = 11'h787 == fractionSum[12:2] ? 10'h3af : _GEN_1926; // @[Multiplier.scala 64:55]
  assign _GEN_1928 = 11'h788 == fractionSum[12:2] ? 10'h3b0 : _GEN_1927; // @[Multiplier.scala 64:55]
  assign _GEN_1929 = 11'h789 == fractionSum[12:2] ? 10'h3b1 : _GEN_1928; // @[Multiplier.scala 64:55]
  assign _GEN_1930 = 11'h78a == fractionSum[12:2] ? 10'h3b1 : _GEN_1929; // @[Multiplier.scala 64:55]
  assign _GEN_1931 = 11'h78b == fractionSum[12:2] ? 10'h3b2 : _GEN_1930; // @[Multiplier.scala 64:55]
  assign _GEN_1932 = 11'h78c == fractionSum[12:2] ? 10'h3b3 : _GEN_1931; // @[Multiplier.scala 64:55]
  assign _GEN_1933 = 11'h78d == fractionSum[12:2] ? 10'h3b3 : _GEN_1932; // @[Multiplier.scala 64:55]
  assign _GEN_1934 = 11'h78e == fractionSum[12:2] ? 10'h3b4 : _GEN_1933; // @[Multiplier.scala 64:55]
  assign _GEN_1935 = 11'h78f == fractionSum[12:2] ? 10'h3b5 : _GEN_1934; // @[Multiplier.scala 64:55]
  assign _GEN_1936 = 11'h790 == fractionSum[12:2] ? 10'h3b5 : _GEN_1935; // @[Multiplier.scala 64:55]
  assign _GEN_1937 = 11'h791 == fractionSum[12:2] ? 10'h3b6 : _GEN_1936; // @[Multiplier.scala 64:55]
  assign _GEN_1938 = 11'h792 == fractionSum[12:2] ? 10'h3b7 : _GEN_1937; // @[Multiplier.scala 64:55]
  assign _GEN_1939 = 11'h793 == fractionSum[12:2] ? 10'h3b7 : _GEN_1938; // @[Multiplier.scala 64:55]
  assign _GEN_1940 = 11'h794 == fractionSum[12:2] ? 10'h3b8 : _GEN_1939; // @[Multiplier.scala 64:55]
  assign _GEN_1941 = 11'h795 == fractionSum[12:2] ? 10'h3b8 : _GEN_1940; // @[Multiplier.scala 64:55]
  assign _GEN_1942 = 11'h796 == fractionSum[12:2] ? 10'h3b9 : _GEN_1941; // @[Multiplier.scala 64:55]
  assign _GEN_1943 = 11'h797 == fractionSum[12:2] ? 10'h3ba : _GEN_1942; // @[Multiplier.scala 64:55]
  assign _GEN_1944 = 11'h798 == fractionSum[12:2] ? 10'h3ba : _GEN_1943; // @[Multiplier.scala 64:55]
  assign _GEN_1945 = 11'h799 == fractionSum[12:2] ? 10'h3bb : _GEN_1944; // @[Multiplier.scala 64:55]
  assign _GEN_1946 = 11'h79a == fractionSum[12:2] ? 10'h3bc : _GEN_1945; // @[Multiplier.scala 64:55]
  assign _GEN_1947 = 11'h79b == fractionSum[12:2] ? 10'h3bc : _GEN_1946; // @[Multiplier.scala 64:55]
  assign _GEN_1948 = 11'h79c == fractionSum[12:2] ? 10'h3bd : _GEN_1947; // @[Multiplier.scala 64:55]
  assign _GEN_1949 = 11'h79d == fractionSum[12:2] ? 10'h3be : _GEN_1948; // @[Multiplier.scala 64:55]
  assign _GEN_1950 = 11'h79e == fractionSum[12:2] ? 10'h3be : _GEN_1949; // @[Multiplier.scala 64:55]
  assign _GEN_1951 = 11'h79f == fractionSum[12:2] ? 10'h3bf : _GEN_1950; // @[Multiplier.scala 64:55]
  assign _GEN_1952 = 11'h7a0 == fractionSum[12:2] ? 10'h3c0 : _GEN_1951; // @[Multiplier.scala 64:55]
  assign _GEN_1953 = 11'h7a1 == fractionSum[12:2] ? 10'h3c0 : _GEN_1952; // @[Multiplier.scala 64:55]
  assign _GEN_1954 = 11'h7a2 == fractionSum[12:2] ? 10'h3c1 : _GEN_1953; // @[Multiplier.scala 64:55]
  assign _GEN_1955 = 11'h7a3 == fractionSum[12:2] ? 10'h3c2 : _GEN_1954; // @[Multiplier.scala 64:55]
  assign _GEN_1956 = 11'h7a4 == fractionSum[12:2] ? 10'h3c2 : _GEN_1955; // @[Multiplier.scala 64:55]
  assign _GEN_1957 = 11'h7a5 == fractionSum[12:2] ? 10'h3c3 : _GEN_1956; // @[Multiplier.scala 64:55]
  assign _GEN_1958 = 11'h7a6 == fractionSum[12:2] ? 10'h3c3 : _GEN_1957; // @[Multiplier.scala 64:55]
  assign _GEN_1959 = 11'h7a7 == fractionSum[12:2] ? 10'h3c4 : _GEN_1958; // @[Multiplier.scala 64:55]
  assign _GEN_1960 = 11'h7a8 == fractionSum[12:2] ? 10'h3c5 : _GEN_1959; // @[Multiplier.scala 64:55]
  assign _GEN_1961 = 11'h7a9 == fractionSum[12:2] ? 10'h3c5 : _GEN_1960; // @[Multiplier.scala 64:55]
  assign _GEN_1962 = 11'h7aa == fractionSum[12:2] ? 10'h3c6 : _GEN_1961; // @[Multiplier.scala 64:55]
  assign _GEN_1963 = 11'h7ab == fractionSum[12:2] ? 10'h3c7 : _GEN_1962; // @[Multiplier.scala 64:55]
  assign _GEN_1964 = 11'h7ac == fractionSum[12:2] ? 10'h3c7 : _GEN_1963; // @[Multiplier.scala 64:55]
  assign _GEN_1965 = 11'h7ad == fractionSum[12:2] ? 10'h3c8 : _GEN_1964; // @[Multiplier.scala 64:55]
  assign _GEN_1966 = 11'h7ae == fractionSum[12:2] ? 10'h3c9 : _GEN_1965; // @[Multiplier.scala 64:55]
  assign _GEN_1967 = 11'h7af == fractionSum[12:2] ? 10'h3c9 : _GEN_1966; // @[Multiplier.scala 64:55]
  assign _GEN_1968 = 11'h7b0 == fractionSum[12:2] ? 10'h3ca : _GEN_1967; // @[Multiplier.scala 64:55]
  assign _GEN_1969 = 11'h7b1 == fractionSum[12:2] ? 10'h3cb : _GEN_1968; // @[Multiplier.scala 64:55]
  assign _GEN_1970 = 11'h7b2 == fractionSum[12:2] ? 10'h3cb : _GEN_1969; // @[Multiplier.scala 64:55]
  assign _GEN_1971 = 11'h7b3 == fractionSum[12:2] ? 10'h3cc : _GEN_1970; // @[Multiplier.scala 64:55]
  assign _GEN_1972 = 11'h7b4 == fractionSum[12:2] ? 10'h3cd : _GEN_1971; // @[Multiplier.scala 64:55]
  assign _GEN_1973 = 11'h7b5 == fractionSum[12:2] ? 10'h3cd : _GEN_1972; // @[Multiplier.scala 64:55]
  assign _GEN_1974 = 11'h7b6 == fractionSum[12:2] ? 10'h3ce : _GEN_1973; // @[Multiplier.scala 64:55]
  assign _GEN_1975 = 11'h7b7 == fractionSum[12:2] ? 10'h3cf : _GEN_1974; // @[Multiplier.scala 64:55]
  assign _GEN_1976 = 11'h7b8 == fractionSum[12:2] ? 10'h3cf : _GEN_1975; // @[Multiplier.scala 64:55]
  assign _GEN_1977 = 11'h7b9 == fractionSum[12:2] ? 10'h3d0 : _GEN_1976; // @[Multiplier.scala 64:55]
  assign _GEN_1978 = 11'h7ba == fractionSum[12:2] ? 10'h3d1 : _GEN_1977; // @[Multiplier.scala 64:55]
  assign _GEN_1979 = 11'h7bb == fractionSum[12:2] ? 10'h3d1 : _GEN_1978; // @[Multiplier.scala 64:55]
  assign _GEN_1980 = 11'h7bc == fractionSum[12:2] ? 10'h3d2 : _GEN_1979; // @[Multiplier.scala 64:55]
  assign _GEN_1981 = 11'h7bd == fractionSum[12:2] ? 10'h3d3 : _GEN_1980; // @[Multiplier.scala 64:55]
  assign _GEN_1982 = 11'h7be == fractionSum[12:2] ? 10'h3d3 : _GEN_1981; // @[Multiplier.scala 64:55]
  assign _GEN_1983 = 11'h7bf == fractionSum[12:2] ? 10'h3d4 : _GEN_1982; // @[Multiplier.scala 64:55]
  assign _GEN_1984 = 11'h7c0 == fractionSum[12:2] ? 10'h3d5 : _GEN_1983; // @[Multiplier.scala 64:55]
  assign _GEN_1985 = 11'h7c1 == fractionSum[12:2] ? 10'h3d5 : _GEN_1984; // @[Multiplier.scala 64:55]
  assign _GEN_1986 = 11'h7c2 == fractionSum[12:2] ? 10'h3d6 : _GEN_1985; // @[Multiplier.scala 64:55]
  assign _GEN_1987 = 11'h7c3 == fractionSum[12:2] ? 10'h3d7 : _GEN_1986; // @[Multiplier.scala 64:55]
  assign _GEN_1988 = 11'h7c4 == fractionSum[12:2] ? 10'h3d7 : _GEN_1987; // @[Multiplier.scala 64:55]
  assign _GEN_1989 = 11'h7c5 == fractionSum[12:2] ? 10'h3d8 : _GEN_1988; // @[Multiplier.scala 64:55]
  assign _GEN_1990 = 11'h7c6 == fractionSum[12:2] ? 10'h3d9 : _GEN_1989; // @[Multiplier.scala 64:55]
  assign _GEN_1991 = 11'h7c7 == fractionSum[12:2] ? 10'h3d9 : _GEN_1990; // @[Multiplier.scala 64:55]
  assign _GEN_1992 = 11'h7c8 == fractionSum[12:2] ? 10'h3da : _GEN_1991; // @[Multiplier.scala 64:55]
  assign _GEN_1993 = 11'h7c9 == fractionSum[12:2] ? 10'h3db : _GEN_1992; // @[Multiplier.scala 64:55]
  assign _GEN_1994 = 11'h7ca == fractionSum[12:2] ? 10'h3db : _GEN_1993; // @[Multiplier.scala 64:55]
  assign _GEN_1995 = 11'h7cb == fractionSum[12:2] ? 10'h3dc : _GEN_1994; // @[Multiplier.scala 64:55]
  assign _GEN_1996 = 11'h7cc == fractionSum[12:2] ? 10'h3dd : _GEN_1995; // @[Multiplier.scala 64:55]
  assign _GEN_1997 = 11'h7cd == fractionSum[12:2] ? 10'h3dd : _GEN_1996; // @[Multiplier.scala 64:55]
  assign _GEN_1998 = 11'h7ce == fractionSum[12:2] ? 10'h3de : _GEN_1997; // @[Multiplier.scala 64:55]
  assign _GEN_1999 = 11'h7cf == fractionSum[12:2] ? 10'h3df : _GEN_1998; // @[Multiplier.scala 64:55]
  assign _GEN_2000 = 11'h7d0 == fractionSum[12:2] ? 10'h3df : _GEN_1999; // @[Multiplier.scala 64:55]
  assign _GEN_2001 = 11'h7d1 == fractionSum[12:2] ? 10'h3e0 : _GEN_2000; // @[Multiplier.scala 64:55]
  assign _GEN_2002 = 11'h7d2 == fractionSum[12:2] ? 10'h3e1 : _GEN_2001; // @[Multiplier.scala 64:55]
  assign _GEN_2003 = 11'h7d3 == fractionSum[12:2] ? 10'h3e1 : _GEN_2002; // @[Multiplier.scala 64:55]
  assign _GEN_2004 = 11'h7d4 == fractionSum[12:2] ? 10'h3e2 : _GEN_2003; // @[Multiplier.scala 64:55]
  assign _GEN_2005 = 11'h7d5 == fractionSum[12:2] ? 10'h3e3 : _GEN_2004; // @[Multiplier.scala 64:55]
  assign _GEN_2006 = 11'h7d6 == fractionSum[12:2] ? 10'h3e3 : _GEN_2005; // @[Multiplier.scala 64:55]
  assign _GEN_2007 = 11'h7d7 == fractionSum[12:2] ? 10'h3e4 : _GEN_2006; // @[Multiplier.scala 64:55]
  assign _GEN_2008 = 11'h7d8 == fractionSum[12:2] ? 10'h3e5 : _GEN_2007; // @[Multiplier.scala 64:55]
  assign _GEN_2009 = 11'h7d9 == fractionSum[12:2] ? 10'h3e5 : _GEN_2008; // @[Multiplier.scala 64:55]
  assign _GEN_2010 = 11'h7da == fractionSum[12:2] ? 10'h3e6 : _GEN_2009; // @[Multiplier.scala 64:55]
  assign _GEN_2011 = 11'h7db == fractionSum[12:2] ? 10'h3e7 : _GEN_2010; // @[Multiplier.scala 64:55]
  assign _GEN_2012 = 11'h7dc == fractionSum[12:2] ? 10'h3e7 : _GEN_2011; // @[Multiplier.scala 64:55]
  assign _GEN_2013 = 11'h7dd == fractionSum[12:2] ? 10'h3e8 : _GEN_2012; // @[Multiplier.scala 64:55]
  assign _GEN_2014 = 11'h7de == fractionSum[12:2] ? 10'h3e9 : _GEN_2013; // @[Multiplier.scala 64:55]
  assign _GEN_2015 = 11'h7df == fractionSum[12:2] ? 10'h3e9 : _GEN_2014; // @[Multiplier.scala 64:55]
  assign _GEN_2016 = 11'h7e0 == fractionSum[12:2] ? 10'h3ea : _GEN_2015; // @[Multiplier.scala 64:55]
  assign _GEN_2017 = 11'h7e1 == fractionSum[12:2] ? 10'h3eb : _GEN_2016; // @[Multiplier.scala 64:55]
  assign _GEN_2018 = 11'h7e2 == fractionSum[12:2] ? 10'h3eb : _GEN_2017; // @[Multiplier.scala 64:55]
  assign _GEN_2019 = 11'h7e3 == fractionSum[12:2] ? 10'h3ec : _GEN_2018; // @[Multiplier.scala 64:55]
  assign _GEN_2020 = 11'h7e4 == fractionSum[12:2] ? 10'h3ed : _GEN_2019; // @[Multiplier.scala 64:55]
  assign _GEN_2021 = 11'h7e5 == fractionSum[12:2] ? 10'h3ed : _GEN_2020; // @[Multiplier.scala 64:55]
  assign _GEN_2022 = 11'h7e6 == fractionSum[12:2] ? 10'h3ee : _GEN_2021; // @[Multiplier.scala 64:55]
  assign _GEN_2023 = 11'h7e7 == fractionSum[12:2] ? 10'h3ef : _GEN_2022; // @[Multiplier.scala 64:55]
  assign _GEN_2024 = 11'h7e8 == fractionSum[12:2] ? 10'h3ef : _GEN_2023; // @[Multiplier.scala 64:55]
  assign _GEN_2025 = 11'h7e9 == fractionSum[12:2] ? 10'h3f0 : _GEN_2024; // @[Multiplier.scala 64:55]
  assign _GEN_2026 = 11'h7ea == fractionSum[12:2] ? 10'h3f1 : _GEN_2025; // @[Multiplier.scala 64:55]
  assign _GEN_2027 = 11'h7eb == fractionSum[12:2] ? 10'h3f2 : _GEN_2026; // @[Multiplier.scala 64:55]
  assign _GEN_2028 = 11'h7ec == fractionSum[12:2] ? 10'h3f2 : _GEN_2027; // @[Multiplier.scala 64:55]
  assign _GEN_2029 = 11'h7ed == fractionSum[12:2] ? 10'h3f3 : _GEN_2028; // @[Multiplier.scala 64:55]
  assign _GEN_2030 = 11'h7ee == fractionSum[12:2] ? 10'h3f4 : _GEN_2029; // @[Multiplier.scala 64:55]
  assign _GEN_2031 = 11'h7ef == fractionSum[12:2] ? 10'h3f4 : _GEN_2030; // @[Multiplier.scala 64:55]
  assign _GEN_2032 = 11'h7f0 == fractionSum[12:2] ? 10'h3f5 : _GEN_2031; // @[Multiplier.scala 64:55]
  assign _GEN_2033 = 11'h7f1 == fractionSum[12:2] ? 10'h3f6 : _GEN_2032; // @[Multiplier.scala 64:55]
  assign _GEN_2034 = 11'h7f2 == fractionSum[12:2] ? 10'h3f6 : _GEN_2033; // @[Multiplier.scala 64:55]
  assign _GEN_2035 = 11'h7f3 == fractionSum[12:2] ? 10'h3f7 : _GEN_2034; // @[Multiplier.scala 64:55]
  assign _GEN_2036 = 11'h7f4 == fractionSum[12:2] ? 10'h3f8 : _GEN_2035; // @[Multiplier.scala 64:55]
  assign _GEN_2037 = 11'h7f5 == fractionSum[12:2] ? 10'h3f8 : _GEN_2036; // @[Multiplier.scala 64:55]
  assign _GEN_2038 = 11'h7f6 == fractionSum[12:2] ? 10'h3f9 : _GEN_2037; // @[Multiplier.scala 64:55]
  assign _GEN_2039 = 11'h7f7 == fractionSum[12:2] ? 10'h3fa : _GEN_2038; // @[Multiplier.scala 64:55]
  assign _GEN_2040 = 11'h7f8 == fractionSum[12:2] ? 10'h3fa : _GEN_2039; // @[Multiplier.scala 64:55]
  assign _GEN_2041 = 11'h7f9 == fractionSum[12:2] ? 10'h3fb : _GEN_2040; // @[Multiplier.scala 64:55]
  assign _GEN_2042 = 11'h7fa == fractionSum[12:2] ? 10'h3fc : _GEN_2041; // @[Multiplier.scala 64:55]
  assign _GEN_2043 = 11'h7fb == fractionSum[12:2] ? 10'h3fd : _GEN_2042; // @[Multiplier.scala 64:55]
  assign _GEN_2044 = 11'h7fc == fractionSum[12:2] ? 10'h3fd : _GEN_2043; // @[Multiplier.scala 64:55]
  assign _GEN_2045 = 11'h7fd == fractionSum[12:2] ? 10'h3fe : _GEN_2044; // @[Multiplier.scala 64:55]
  assign _GEN_2046 = 11'h7fe == fractionSum[12:2] ? 10'h3ff : _GEN_2045; // @[Multiplier.scala 64:55]
  assign _GEN_2047 = 11'h7ff == fractionSum[12:2] ? 10'h3ff : _GEN_2046; // @[Multiplier.scala 64:55]
  assign _T_10 = _GEN_2047 >> _T_9; // @[Multiplier.scala 64:55]
  assign _T_11 = $signed(_T_4) - 8'sh8; // @[Multiplier.scala 64:100]
  assign _GEN_2048 = {{511'd0}, _GEN_2047}; // @[Multiplier.scala 64:91]
  assign _T_12 = _GEN_2048 << _T_11; // @[Multiplier.scala 64:91]
  assign _T_13 = io_A_zero | io_B_zero; // @[Multiplier.scala 66:34]
  assign _T_16 = 6'sh0 - 6'sh18; // @[Multiplier.scala 66:57]
  assign _GEN_2049 = {{3{_T_16[5]}},_T_16}; // @[Multiplier.scala 66:55]
  assign _T_17 = $signed(shift) < $signed(_GEN_2049); // @[Multiplier.scala 66:55]
  assign _T_19 = io_A_nan | io_B_nan; // @[Multiplier.scala 67:32]
  assign _T_20 = $signed(shift) >= 9'sh77; // @[Multiplier.scala 67:52]
  assign _T_22 = io_out_zero | io_out_nan; // @[Multiplier.scala 68:42]
  assign _T_23 = io_A_sign ^ io_B_sign; // @[Multiplier.scala 68:76]
  assign _T_25 = _T_5 ? {{511'd0}, _T_10} : _T_12; // @[Multiplier.scala 68:105]
  assign _T_28 = 521'sh0 - $signed(_T_25); // @[Multiplier.scala 68:97]
  assign _T_30 = _T_23 ? $signed(_T_28) : $signed(_T_25); // @[Multiplier.scala 68:64]
  assign _T_31 = _T_22 ? $signed(521'sh0) : $signed(_T_30); // @[Multiplier.scala 68:29]
  assign io_out_zero = _T_13 | _T_17; // @[Multiplier.scala 66:21]
  assign io_out_nan = _T_19 | _T_20; // @[Multiplier.scala 67:20]
  assign io_out_number = _T_31[128:0]; // @[Multiplier.scala 68:23]
endmodule
module logMultiplierMAC(
  input          io_A_zero,
  input          io_A_nan,
  input          io_A_sign,
  input  [5:0]   io_A_exponent,
  input  [12:0]  io_A_fraction,
  input          io_B_zero,
  input          io_B_nan,
  input          io_B_sign,
  input  [5:0]   io_B_exponent,
  input  [12:0]  io_B_fraction,
  input          io_C_zero,
  input          io_C_nan,
  input  [128:0] io_C_number,
  output         io_out_zero,
  output         io_out_nan,
  output [128:0] io_out_number
);
  wire  multiplier_io_A_zero; // @[Multiplier.scala 79:32]
  wire  multiplier_io_A_nan; // @[Multiplier.scala 79:32]
  wire  multiplier_io_A_sign; // @[Multiplier.scala 79:32]
  wire [5:0] multiplier_io_A_exponent; // @[Multiplier.scala 79:32]
  wire [12:0] multiplier_io_A_fraction; // @[Multiplier.scala 79:32]
  wire  multiplier_io_B_zero; // @[Multiplier.scala 79:32]
  wire  multiplier_io_B_nan; // @[Multiplier.scala 79:32]
  wire  multiplier_io_B_sign; // @[Multiplier.scala 79:32]
  wire [5:0] multiplier_io_B_exponent; // @[Multiplier.scala 79:32]
  wire [12:0] multiplier_io_B_fraction; // @[Multiplier.scala 79:32]
  wire  multiplier_io_out_zero; // @[Multiplier.scala 79:32]
  wire  multiplier_io_out_nan; // @[Multiplier.scala 79:32]
  wire [128:0] multiplier_io_out_number; // @[Multiplier.scala 79:32]
  wire [128:0] sum; // @[Multiplier.scala 82:44]
  wire  _T_2; // @[Multiplier.scala 83:48]
  wire  _T_5; // @[Multiplier.scala 83:99]
  wire  _T_8; // @[Multiplier.scala 83:151]
  wire  _T_10; // @[Multiplier.scala 83:228]
  wire  _T_11; // @[Multiplier.scala 83:198]
  wire  _T_13; // @[Multiplier.scala 84:45]
  wire  _T_18; // @[Multiplier.scala 84:184]
  wire  _T_19; // @[Multiplier.scala 84:146]
  wire  _T_22; // @[Multiplier.scala 84:193]
  logMultiplier multiplier ( // @[Multiplier.scala 79:32]
    .io_A_zero(multiplier_io_A_zero),
    .io_A_nan(multiplier_io_A_nan),
    .io_A_sign(multiplier_io_A_sign),
    .io_A_exponent(multiplier_io_A_exponent),
    .io_A_fraction(multiplier_io_A_fraction),
    .io_B_zero(multiplier_io_B_zero),
    .io_B_nan(multiplier_io_B_nan),
    .io_B_sign(multiplier_io_B_sign),
    .io_B_exponent(multiplier_io_B_exponent),
    .io_B_fraction(multiplier_io_B_fraction),
    .io_out_zero(multiplier_io_out_zero),
    .io_out_nan(multiplier_io_out_nan),
    .io_out_number(multiplier_io_out_number)
  );
  assign sum = $signed(multiplier_io_out_number) + $signed(io_C_number); // @[Multiplier.scala 82:44]
  assign _T_2 = multiplier_io_out_zero & io_C_zero; // @[Multiplier.scala 83:48]
  assign _T_5 = io_C_number[128] == multiplier_io_out_number[128]; // @[Multiplier.scala 83:99]
  assign _T_8 = _T_5 & io_C_number[128]; // @[Multiplier.scala 83:151]
  assign _T_10 = ~sum[128]; // @[Multiplier.scala 83:228]
  assign _T_11 = _T_8 & _T_10; // @[Multiplier.scala 83:198]
  assign _T_13 = multiplier_io_out_nan | io_C_nan; // @[Multiplier.scala 84:45]
  assign _T_18 = ~io_C_number[128]; // @[Multiplier.scala 84:184]
  assign _T_19 = _T_5 & _T_18; // @[Multiplier.scala 84:146]
  assign _T_22 = _T_19 & sum[128]; // @[Multiplier.scala 84:193]
  assign io_out_zero = _T_2 | _T_11; // @[Multiplier.scala 83:21]
  assign io_out_nan = _T_13 | _T_22; // @[Multiplier.scala 84:20]
  assign io_out_number = $signed(multiplier_io_out_number) + $signed(io_C_number); // @[Multiplier.scala 85:23]
  assign multiplier_io_A_zero = io_A_zero; // @[Multiplier.scala 80:25]
  assign multiplier_io_A_nan = io_A_nan; // @[Multiplier.scala 80:25]
  assign multiplier_io_A_sign = io_A_sign; // @[Multiplier.scala 80:25]
  assign multiplier_io_A_exponent = io_A_exponent; // @[Multiplier.scala 80:25]
  assign multiplier_io_A_fraction = io_A_fraction; // @[Multiplier.scala 80:25]
  assign multiplier_io_B_zero = io_B_zero; // @[Multiplier.scala 81:25]
  assign multiplier_io_B_nan = io_B_nan; // @[Multiplier.scala 81:25]
  assign multiplier_io_B_sign = io_B_sign; // @[Multiplier.scala 81:25]
  assign multiplier_io_B_exponent = io_B_exponent; // @[Multiplier.scala 81:25]
  assign multiplier_io_B_fraction = io_B_fraction; // @[Multiplier.scala 81:25]
endmodule
module logTile(
  input          clock,
  input          io_A_in_zero,
  input          io_A_in_nan,
  input          io_A_in_sign,
  input  [5:0]   io_A_in_exponent,
  input  [12:0]  io_A_in_fraction,
  input          io_B_in_zero,
  input          io_B_in_nan,
  input          io_B_in_sign,
  input  [5:0]   io_B_in_exponent,
  input  [12:0]  io_B_in_fraction,
  input          io_C_in_zero,
  input          io_C_in_nan,
  input  [128:0] io_C_in_number,
  input          io_prop_in,
  output         io_A_out_zero,
  output         io_A_out_nan,
  output         io_A_out_sign,
  output [5:0]   io_A_out_exponent,
  output [12:0]  io_A_out_fraction,
  output         io_B_out_zero,
  output         io_B_out_nan,
  output         io_B_out_sign,
  output [5:0]   io_B_out_exponent,
  output [12:0]  io_B_out_fraction,
  output         io_C_out_zero,
  output         io_C_out_nan,
  output [128:0] io_C_out_number,
  output         io_prop_out
);
  wire  mac_io_A_zero; // @[Tile.scala 65:33]
  wire  mac_io_A_nan; // @[Tile.scala 65:33]
  wire  mac_io_A_sign; // @[Tile.scala 65:33]
  wire [5:0] mac_io_A_exponent; // @[Tile.scala 65:33]
  wire [12:0] mac_io_A_fraction; // @[Tile.scala 65:33]
  wire  mac_io_B_zero; // @[Tile.scala 65:33]
  wire  mac_io_B_nan; // @[Tile.scala 65:33]
  wire  mac_io_B_sign; // @[Tile.scala 65:33]
  wire [5:0] mac_io_B_exponent; // @[Tile.scala 65:33]
  wire [12:0] mac_io_B_fraction; // @[Tile.scala 65:33]
  wire  mac_io_C_zero; // @[Tile.scala 65:33]
  wire  mac_io_C_nan; // @[Tile.scala 65:33]
  wire [128:0] mac_io_C_number; // @[Tile.scala 65:33]
  wire  mac_io_out_zero; // @[Tile.scala 65:33]
  wire  mac_io_out_nan; // @[Tile.scala 65:33]
  wire [128:0] mac_io_out_number; // @[Tile.scala 65:33]
  wire  _T; // @[Tile.scala 58:45]
  reg  A0_zero; // @[Reg.scala 15:16]
  reg [31:0] _RAND_0;
  reg  A0_nan; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1;
  reg  A0_sign; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2;
  reg [5:0] A0_exponent; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3;
  reg [12:0] A0_fraction; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4;
  reg  A1_zero; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5;
  reg  A1_nan; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6;
  reg  A1_sign; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7;
  reg [5:0] A1_exponent; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8;
  reg [12:0] A1_fraction; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9;
  reg  A_zero; // @[Tile.scala 61:32]
  reg [31:0] _RAND_10;
  reg  A_nan; // @[Tile.scala 61:32]
  reg [31:0] _RAND_11;
  reg  A_sign; // @[Tile.scala 61:32]
  reg [31:0] _RAND_12;
  reg [5:0] A_exponent; // @[Tile.scala 61:32]
  reg [31:0] _RAND_13;
  reg [12:0] A_fraction; // @[Tile.scala 61:32]
  reg [31:0] _RAND_14;
  reg  B_zero; // @[Tile.scala 62:32]
  reg [31:0] _RAND_15;
  reg  B_nan; // @[Tile.scala 62:32]
  reg [31:0] _RAND_16;
  reg  B_sign; // @[Tile.scala 62:32]
  reg [31:0] _RAND_17;
  reg [5:0] B_exponent; // @[Tile.scala 62:32]
  reg [31:0] _RAND_18;
  reg [12:0] B_fraction; // @[Tile.scala 62:32]
  reg [31:0] _RAND_19;
  reg  prop; // @[Tile.scala 63:35]
  reg [31:0] _RAND_20;
  reg  C_zero; // @[Tile.scala 70:32]
  reg [31:0] _RAND_21;
  reg  C_nan; // @[Tile.scala 70:32]
  reg [31:0] _RAND_22;
  reg [128:0] C_number; // @[Tile.scala 70:32]
  reg [159:0] _RAND_23;
  logMultiplierMAC mac ( // @[Tile.scala 65:33]
    .io_A_zero(mac_io_A_zero),
    .io_A_nan(mac_io_A_nan),
    .io_A_sign(mac_io_A_sign),
    .io_A_exponent(mac_io_A_exponent),
    .io_A_fraction(mac_io_A_fraction),
    .io_B_zero(mac_io_B_zero),
    .io_B_nan(mac_io_B_nan),
    .io_B_sign(mac_io_B_sign),
    .io_B_exponent(mac_io_B_exponent),
    .io_B_fraction(mac_io_B_fraction),
    .io_C_zero(mac_io_C_zero),
    .io_C_nan(mac_io_C_nan),
    .io_C_number(mac_io_C_number),
    .io_out_zero(mac_io_out_zero),
    .io_out_nan(mac_io_out_nan),
    .io_out_number(mac_io_out_number)
  );
  assign _T = ~io_prop_in; // @[Tile.scala 58:45]
  assign io_A_out_zero = A_zero; // @[Tile.scala 72:26]
  assign io_A_out_nan = A_nan; // @[Tile.scala 72:26]
  assign io_A_out_sign = A_sign; // @[Tile.scala 72:26]
  assign io_A_out_exponent = A_exponent; // @[Tile.scala 72:26]
  assign io_A_out_fraction = A_fraction; // @[Tile.scala 72:26]
  assign io_B_out_zero = B_zero; // @[Tile.scala 73:26]
  assign io_B_out_nan = B_nan; // @[Tile.scala 73:26]
  assign io_B_out_sign = B_sign; // @[Tile.scala 73:26]
  assign io_B_out_exponent = B_exponent; // @[Tile.scala 73:26]
  assign io_B_out_fraction = B_fraction; // @[Tile.scala 73:26]
  assign io_C_out_zero = C_zero; // @[Tile.scala 74:26]
  assign io_C_out_nan = C_nan; // @[Tile.scala 74:26]
  assign io_C_out_number = C_number; // @[Tile.scala 74:26]
  assign io_prop_out = prop; // @[Tile.scala 75:29]
  assign mac_io_A_zero = io_prop_in ? A0_zero : A1_zero; // @[Tile.scala 66:26]
  assign mac_io_A_nan = io_prop_in ? A0_nan : A1_nan; // @[Tile.scala 66:26]
  assign mac_io_A_sign = io_prop_in ? A0_sign : A1_sign; // @[Tile.scala 66:26]
  assign mac_io_A_exponent = io_prop_in ? $signed(A0_exponent) : $signed(A1_exponent); // @[Tile.scala 66:26]
  assign mac_io_A_fraction = io_prop_in ? A0_fraction : A1_fraction; // @[Tile.scala 66:26]
  assign mac_io_B_zero = io_B_in_zero; // @[Tile.scala 67:26]
  assign mac_io_B_nan = io_B_in_nan; // @[Tile.scala 67:26]
  assign mac_io_B_sign = io_B_in_sign; // @[Tile.scala 67:26]
  assign mac_io_B_exponent = io_B_in_exponent; // @[Tile.scala 67:26]
  assign mac_io_B_fraction = io_B_in_fraction; // @[Tile.scala 67:26]
  assign mac_io_C_zero = io_C_in_zero; // @[Tile.scala 68:26]
  assign mac_io_C_nan = io_C_in_nan; // @[Tile.scala 68:26]
  assign mac_io_C_number = io_C_in_number; // @[Tile.scala 68:26]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  A0_zero = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  A0_nan = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  A0_sign = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  A0_exponent = _RAND_3[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  A0_fraction = _RAND_4[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  A1_zero = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  A1_nan = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  A1_sign = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  A1_exponent = _RAND_8[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  A1_fraction = _RAND_9[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  A_zero = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  A_nan = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  A_sign = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  A_exponent = _RAND_13[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  A_fraction = _RAND_14[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  B_zero = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  B_nan = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  B_sign = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  B_exponent = _RAND_18[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  B_fraction = _RAND_19[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  prop = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  C_zero = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  C_nan = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {5{`RANDOM}};
  C_number = _RAND_23[128:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (_T) begin
      A0_zero <= io_A_in_zero;
    end
    if (_T) begin
      A0_nan <= io_A_in_nan;
    end
    if (_T) begin
      A0_sign <= io_A_in_sign;
    end
    if (_T) begin
      A0_exponent <= io_A_in_exponent;
    end
    if (_T) begin
      A0_fraction <= io_A_in_fraction;
    end
    if (io_prop_in) begin
      A1_zero <= io_A_in_zero;
    end
    if (io_prop_in) begin
      A1_nan <= io_A_in_nan;
    end
    if (io_prop_in) begin
      A1_sign <= io_A_in_sign;
    end
    if (io_prop_in) begin
      A1_exponent <= io_A_in_exponent;
    end
    if (io_prop_in) begin
      A1_fraction <= io_A_in_fraction;
    end
    if (io_prop_in) begin
      A_zero <= A1_zero;
    end else begin
      A_zero <= A0_zero;
    end
    if (io_prop_in) begin
      A_nan <= A1_nan;
    end else begin
      A_nan <= A0_nan;
    end
    if (io_prop_in) begin
      A_sign <= A1_sign;
    end else begin
      A_sign <= A0_sign;
    end
    if (io_prop_in) begin
      A_exponent <= A1_exponent;
    end else begin
      A_exponent <= A0_exponent;
    end
    if (io_prop_in) begin
      A_fraction <= A1_fraction;
    end else begin
      A_fraction <= A0_fraction;
    end
    B_zero <= io_B_in_zero;
    B_nan <= io_B_in_nan;
    B_sign <= io_B_in_sign;
    B_exponent <= io_B_in_exponent;
    B_fraction <= io_B_in_fraction;
    prop <= io_prop_in;
    C_zero <= mac_io_out_zero;
    C_nan <= mac_io_out_nan;
    C_number <= mac_io_out_number;
  end
endmodule
module toPositUnpacked(
  input  [15:0] io_in,
  output        io_out_zero,
  output        io_out_nan,
  output        io_out_sign,
  output [5:0]  io_out_exponent,
  output [12:0] io_out_fraction
);
  wire [14:0] _T_2; // @[Bitwise.scala 71:12]
  wire [14:0] _T_3; // @[Conversion.scala 20:43]
  wire [14:0] _GEN_0; // @[Conversion.scala 20:78]
  wire [14:0] others; // @[Conversion.scala 20:78]
  wire [14:0] _T_7; // @[Conversion.scala 21:77]
  wire [7:0] _T_12; // @[Bitwise.scala 102:31]
  wire [7:0] _T_14; // @[Bitwise.scala 102:65]
  wire [7:0] _T_16; // @[Bitwise.scala 102:75]
  wire [7:0] _T_17; // @[Bitwise.scala 102:39]
  wire [7:0] _GEN_1; // @[Bitwise.scala 102:31]
  wire [7:0] _T_22; // @[Bitwise.scala 102:31]
  wire [7:0] _T_24; // @[Bitwise.scala 102:65]
  wire [7:0] _T_26; // @[Bitwise.scala 102:75]
  wire [7:0] _T_27; // @[Bitwise.scala 102:39]
  wire [7:0] _GEN_2; // @[Bitwise.scala 102:31]
  wire [7:0] _T_32; // @[Bitwise.scala 102:31]
  wire [7:0] _T_34; // @[Bitwise.scala 102:65]
  wire [7:0] _T_36; // @[Bitwise.scala 102:75]
  wire [7:0] _T_37; // @[Bitwise.scala 102:39]
  wire [14:0] _T_57; // @[Cat.scala 29:58]
  wire [3:0] _T_73; // @[Mux.scala 47:69]
  wire [3:0] _T_74; // @[Mux.scala 47:69]
  wire [3:0] _T_75; // @[Mux.scala 47:69]
  wire [3:0] _T_76; // @[Mux.scala 47:69]
  wire [3:0] _T_77; // @[Mux.scala 47:69]
  wire [3:0] _T_78; // @[Mux.scala 47:69]
  wire [3:0] _T_79; // @[Mux.scala 47:69]
  wire [3:0] _T_80; // @[Mux.scala 47:69]
  wire [3:0] _T_81; // @[Mux.scala 47:69]
  wire [3:0] _T_82; // @[Mux.scala 47:69]
  wire [3:0] _T_83; // @[Mux.scala 47:69]
  wire [3:0] _T_84; // @[Mux.scala 47:69]
  wire [3:0] _T_85; // @[Mux.scala 47:69]
  wire [3:0] _T_86; // @[Mux.scala 47:69]
  wire [7:0] _T_91; // @[Bitwise.scala 102:31]
  wire [7:0] _T_93; // @[Bitwise.scala 102:65]
  wire [7:0] _T_95; // @[Bitwise.scala 102:75]
  wire [7:0] _T_96; // @[Bitwise.scala 102:39]
  wire [7:0] _GEN_3; // @[Bitwise.scala 102:31]
  wire [7:0] _T_101; // @[Bitwise.scala 102:31]
  wire [7:0] _T_103; // @[Bitwise.scala 102:65]
  wire [7:0] _T_105; // @[Bitwise.scala 102:75]
  wire [7:0] _T_106; // @[Bitwise.scala 102:39]
  wire [7:0] _GEN_4; // @[Bitwise.scala 102:31]
  wire [7:0] _T_111; // @[Bitwise.scala 102:31]
  wire [7:0] _T_113; // @[Bitwise.scala 102:65]
  wire [7:0] _T_115; // @[Bitwise.scala 102:75]
  wire [7:0] _T_116; // @[Bitwise.scala 102:39]
  wire [14:0] _T_136; // @[Cat.scala 29:58]
  wire [3:0] _T_152; // @[Mux.scala 47:69]
  wire [3:0] _T_153; // @[Mux.scala 47:69]
  wire [3:0] _T_154; // @[Mux.scala 47:69]
  wire [3:0] _T_155; // @[Mux.scala 47:69]
  wire [3:0] _T_156; // @[Mux.scala 47:69]
  wire [3:0] _T_157; // @[Mux.scala 47:69]
  wire [3:0] _T_158; // @[Mux.scala 47:69]
  wire [3:0] _T_159; // @[Mux.scala 47:69]
  wire [3:0] _T_160; // @[Mux.scala 47:69]
  wire [3:0] _T_161; // @[Mux.scala 47:69]
  wire [3:0] _T_162; // @[Mux.scala 47:69]
  wire [3:0] _T_163; // @[Mux.scala 47:69]
  wire [3:0] _T_164; // @[Mux.scala 47:69]
  wire [3:0] _T_165; // @[Mux.scala 47:69]
  wire [3:0] _T_166; // @[Conversion.scala 21:23]
  wire  _T_167; // @[Conversion.scala 21:132]
  wire  _T_168; // @[Conversion.scala 21:147]
  wire  _T_169; // @[Conversion.scala 21:139]
  wire  _T_170; // @[Conversion.scala 21:137]
  wire [3:0] _GEN_5; // @[Conversion.scala 21:122]
  wire [3:0] _T_172; // @[Conversion.scala 21:122]
  wire [4:0] leading; // @[Conversion.scala 14:27 Conversion.scala 21:17]
  wire [4:0] _T_174; // @[Conversion.scala 22:60]
  wire [4:0] _T_177; // @[Conversion.scala 22:67]
  wire [4:0] _T_181; // @[Conversion.scala 22:74]
  wire [4:0] _T_182; // @[Conversion.scala 22:22]
  wire [4:0] _T_184; // @[Conversion.scala 23:48]
  wire [45:0] _GEN_6; // @[Conversion.scala 23:36]
  wire [45:0] _T_185; // @[Conversion.scala 23:36]
  wire [12:0] exponentFraction; // @[Conversion.scala 16:36 Conversion.scala 23:26]
  wire  exponent; // @[Conversion.scala 24:37]
  wire  _T_190; // @[Conversion.scala 27:24]
  wire  _T_192; // @[Conversion.scala 27:71]
  wire  _T_193; // @[Conversion.scala 27:47]
  wire [5:0] regime; // @[Conversion.scala 15:26 Conversion.scala 22:16]
  wire [6:0] _T_201; // @[Conversion.scala 30:36]
  wire [1:0] _T_202; // @[Conversion.scala 30:99]
  wire [6:0] _GEN_7; // @[Conversion.scala 30:88]
  wire [6:0] _T_205; // @[Conversion.scala 30:88]
  assign _T_2 = io_out_sign ? 15'h7fff : 15'h0; // @[Bitwise.scala 71:12]
  assign _T_3 = io_in[14:0] ^ _T_2; // @[Conversion.scala 20:43]
  assign _GEN_0 = {{14'd0}, io_out_sign}; // @[Conversion.scala 20:78]
  assign others = _T_3 + _GEN_0; // @[Conversion.scala 20:78]
  assign _T_7 = ~others; // @[Conversion.scala 21:77]
  assign _T_12 = {{4'd0}, _T_7[7:4]}; // @[Bitwise.scala 102:31]
  assign _T_14 = {_T_7[3:0], 4'h0}; // @[Bitwise.scala 102:65]
  assign _T_16 = _T_14 & 8'hf0; // @[Bitwise.scala 102:75]
  assign _T_17 = _T_12 | _T_16; // @[Bitwise.scala 102:39]
  assign _GEN_1 = {{2'd0}, _T_17[7:2]}; // @[Bitwise.scala 102:31]
  assign _T_22 = _GEN_1 & 8'h33; // @[Bitwise.scala 102:31]
  assign _T_24 = {_T_17[5:0], 2'h0}; // @[Bitwise.scala 102:65]
  assign _T_26 = _T_24 & 8'hcc; // @[Bitwise.scala 102:75]
  assign _T_27 = _T_22 | _T_26; // @[Bitwise.scala 102:39]
  assign _GEN_2 = {{1'd0}, _T_27[7:1]}; // @[Bitwise.scala 102:31]
  assign _T_32 = _GEN_2 & 8'h55; // @[Bitwise.scala 102:31]
  assign _T_34 = {_T_27[6:0], 1'h0}; // @[Bitwise.scala 102:65]
  assign _T_36 = _T_34 & 8'haa; // @[Bitwise.scala 102:75]
  assign _T_37 = _T_32 | _T_36; // @[Bitwise.scala 102:39]
  assign _T_57 = {_T_37,_T_7[8],_T_7[9],_T_7[10],_T_7[11],_T_7[12],_T_7[13],_T_7[14]}; // @[Cat.scala 29:58]
  assign _T_73 = _T_57[13] ? 4'hd : 4'he; // @[Mux.scala 47:69]
  assign _T_74 = _T_57[12] ? 4'hc : _T_73; // @[Mux.scala 47:69]
  assign _T_75 = _T_57[11] ? 4'hb : _T_74; // @[Mux.scala 47:69]
  assign _T_76 = _T_57[10] ? 4'ha : _T_75; // @[Mux.scala 47:69]
  assign _T_77 = _T_57[9] ? 4'h9 : _T_76; // @[Mux.scala 47:69]
  assign _T_78 = _T_57[8] ? 4'h8 : _T_77; // @[Mux.scala 47:69]
  assign _T_79 = _T_57[7] ? 4'h7 : _T_78; // @[Mux.scala 47:69]
  assign _T_80 = _T_57[6] ? 4'h6 : _T_79; // @[Mux.scala 47:69]
  assign _T_81 = _T_57[5] ? 4'h5 : _T_80; // @[Mux.scala 47:69]
  assign _T_82 = _T_57[4] ? 4'h4 : _T_81; // @[Mux.scala 47:69]
  assign _T_83 = _T_57[3] ? 4'h3 : _T_82; // @[Mux.scala 47:69]
  assign _T_84 = _T_57[2] ? 4'h2 : _T_83; // @[Mux.scala 47:69]
  assign _T_85 = _T_57[1] ? 4'h1 : _T_84; // @[Mux.scala 47:69]
  assign _T_86 = _T_57[0] ? 4'h0 : _T_85; // @[Mux.scala 47:69]
  assign _T_91 = {{4'd0}, others[7:4]}; // @[Bitwise.scala 102:31]
  assign _T_93 = {others[3:0], 4'h0}; // @[Bitwise.scala 102:65]
  assign _T_95 = _T_93 & 8'hf0; // @[Bitwise.scala 102:75]
  assign _T_96 = _T_91 | _T_95; // @[Bitwise.scala 102:39]
  assign _GEN_3 = {{2'd0}, _T_96[7:2]}; // @[Bitwise.scala 102:31]
  assign _T_101 = _GEN_3 & 8'h33; // @[Bitwise.scala 102:31]
  assign _T_103 = {_T_96[5:0], 2'h0}; // @[Bitwise.scala 102:65]
  assign _T_105 = _T_103 & 8'hcc; // @[Bitwise.scala 102:75]
  assign _T_106 = _T_101 | _T_105; // @[Bitwise.scala 102:39]
  assign _GEN_4 = {{1'd0}, _T_106[7:1]}; // @[Bitwise.scala 102:31]
  assign _T_111 = _GEN_4 & 8'h55; // @[Bitwise.scala 102:31]
  assign _T_113 = {_T_106[6:0], 1'h0}; // @[Bitwise.scala 102:65]
  assign _T_115 = _T_113 & 8'haa; // @[Bitwise.scala 102:75]
  assign _T_116 = _T_111 | _T_115; // @[Bitwise.scala 102:39]
  assign _T_136 = {_T_116,others[8],others[9],others[10],others[11],others[12],others[13],others[14]}; // @[Cat.scala 29:58]
  assign _T_152 = _T_136[13] ? 4'hd : 4'he; // @[Mux.scala 47:69]
  assign _T_153 = _T_136[12] ? 4'hc : _T_152; // @[Mux.scala 47:69]
  assign _T_154 = _T_136[11] ? 4'hb : _T_153; // @[Mux.scala 47:69]
  assign _T_155 = _T_136[10] ? 4'ha : _T_154; // @[Mux.scala 47:69]
  assign _T_156 = _T_136[9] ? 4'h9 : _T_155; // @[Mux.scala 47:69]
  assign _T_157 = _T_136[8] ? 4'h8 : _T_156; // @[Mux.scala 47:69]
  assign _T_158 = _T_136[7] ? 4'h7 : _T_157; // @[Mux.scala 47:69]
  assign _T_159 = _T_136[6] ? 4'h6 : _T_158; // @[Mux.scala 47:69]
  assign _T_160 = _T_136[5] ? 4'h5 : _T_159; // @[Mux.scala 47:69]
  assign _T_161 = _T_136[4] ? 4'h4 : _T_160; // @[Mux.scala 47:69]
  assign _T_162 = _T_136[3] ? 4'h3 : _T_161; // @[Mux.scala 47:69]
  assign _T_163 = _T_136[2] ? 4'h2 : _T_162; // @[Mux.scala 47:69]
  assign _T_164 = _T_136[1] ? 4'h1 : _T_163; // @[Mux.scala 47:69]
  assign _T_165 = _T_136[0] ? 4'h0 : _T_164; // @[Mux.scala 47:69]
  assign _T_166 = others[14] ? _T_86 : _T_165; // @[Conversion.scala 21:23]
  assign _T_167 = others == 15'h7fff; // @[Conversion.scala 21:132]
  assign _T_168 = others != 15'h0; // @[Conversion.scala 21:147]
  assign _T_169 = ~_T_168; // @[Conversion.scala 21:139]
  assign _T_170 = _T_167 | _T_169; // @[Conversion.scala 21:137]
  assign _GEN_5 = {{3'd0}, _T_170}; // @[Conversion.scala 21:122]
  assign _T_172 = _T_166 + _GEN_5; // @[Conversion.scala 21:122]
  assign leading = {{1'd0}, _T_172}; // @[Conversion.scala 14:27 Conversion.scala 21:17]
  assign _T_174 = {{1'd0}, _T_172}; // @[Conversion.scala 22:60]
  assign _T_177 = $signed(_T_174) - 5'sh1; // @[Conversion.scala 22:67]
  assign _T_181 = 5'sh0 - $signed(_T_174); // @[Conversion.scala 22:74]
  assign _T_182 = others[14] ? $signed(_T_177) : $signed(_T_181); // @[Conversion.scala 22:22]
  assign _T_184 = leading - 5'h1; // @[Conversion.scala 23:48]
  assign _GEN_6 = {{31'd0}, others}; // @[Conversion.scala 23:36]
  assign _T_185 = _GEN_6 << _T_184; // @[Conversion.scala 23:36]
  assign exponentFraction = _T_185[12:0]; // @[Conversion.scala 16:36 Conversion.scala 23:26]
  assign exponent = exponentFraction[12]; // @[Conversion.scala 24:37]
  assign _T_190 = ~io_in[15]; // @[Conversion.scala 27:24]
  assign _T_192 = io_in[14:0] != 15'h0; // @[Conversion.scala 27:71]
  assign _T_193 = ~_T_192; // @[Conversion.scala 27:47]
  assign regime = {{1{_T_182[4]}},_T_182}; // @[Conversion.scala 15:26 Conversion.scala 22:16]
  assign _T_201 = {$signed(regime), 1'h0}; // @[Conversion.scala 30:36]
  assign _T_202 = {1'b0,$signed(exponent)}; // @[Conversion.scala 30:99]
  assign _GEN_7 = {{5{_T_202[1]}},_T_202}; // @[Conversion.scala 30:88]
  assign _T_205 = $signed(_T_201) + $signed(_GEN_7); // @[Conversion.scala 30:88]
  assign io_out_zero = _T_190 & _T_193; // @[Conversion.scala 27:21]
  assign io_out_nan = io_in[15] & _T_193; // @[Conversion.scala 28:20]
  assign io_out_sign = io_in[15]; // @[Conversion.scala 29:21]
  assign io_out_exponent = _T_205[5:0]; // @[Conversion.scala 30:25]
  assign io_out_fraction = {1'h1,exponentFraction[11:0]}; // @[Conversion.scala 31:25]
endmodule
module logPositArray(
  input          clock,
  input          reset,
  input  [15:0]  io_A_in_0,
  input  [15:0]  io_A_in_1,
  input  [15:0]  io_A_in_2,
  input  [15:0]  io_A_in_3,
  input  [15:0]  io_B_in_0,
  input  [15:0]  io_B_in_1,
  input  [15:0]  io_B_in_2,
  input  [15:0]  io_B_in_3,
  input          io_C_in_0_zero,
  input          io_C_in_0_nan,
  input  [128:0] io_C_in_0_number,
  input          io_C_in_1_zero,
  input          io_C_in_1_nan,
  input  [128:0] io_C_in_1_number,
  input          io_C_in_2_zero,
  input          io_C_in_2_nan,
  input  [128:0] io_C_in_2_number,
  input          io_C_in_3_zero,
  input          io_C_in_3_nan,
  input  [128:0] io_C_in_3_number,
  input          io_prop_in_0,
  input          io_prop_in_1,
  input          io_prop_in_2,
  input          io_prop_in_3,
  output         io_C_out_0_zero,
  output         io_C_out_0_nan,
  output [128:0] io_C_out_0_number,
  output         io_C_out_1_zero,
  output         io_C_out_1_nan,
  output [128:0] io_C_out_1_number,
  output         io_C_out_2_zero,
  output         io_C_out_2_nan,
  output [128:0] io_C_out_2_number,
  output         io_C_out_3_zero,
  output         io_C_out_3_nan,
  output [128:0] io_C_out_3_number
);
  wire  array_0_0_clock; // @[Array.scala 95:75]
  wire  array_0_0_io_A_in_zero; // @[Array.scala 95:75]
  wire  array_0_0_io_A_in_nan; // @[Array.scala 95:75]
  wire  array_0_0_io_A_in_sign; // @[Array.scala 95:75]
  wire [5:0] array_0_0_io_A_in_exponent; // @[Array.scala 95:75]
  wire [12:0] array_0_0_io_A_in_fraction; // @[Array.scala 95:75]
  wire  array_0_0_io_B_in_zero; // @[Array.scala 95:75]
  wire  array_0_0_io_B_in_nan; // @[Array.scala 95:75]
  wire  array_0_0_io_B_in_sign; // @[Array.scala 95:75]
  wire [5:0] array_0_0_io_B_in_exponent; // @[Array.scala 95:75]
  wire [12:0] array_0_0_io_B_in_fraction; // @[Array.scala 95:75]
  wire  array_0_0_io_C_in_zero; // @[Array.scala 95:75]
  wire  array_0_0_io_C_in_nan; // @[Array.scala 95:75]
  wire [128:0] array_0_0_io_C_in_number; // @[Array.scala 95:75]
  wire  array_0_0_io_prop_in; // @[Array.scala 95:75]
  wire  array_0_0_io_A_out_zero; // @[Array.scala 95:75]
  wire  array_0_0_io_A_out_nan; // @[Array.scala 95:75]
  wire  array_0_0_io_A_out_sign; // @[Array.scala 95:75]
  wire [5:0] array_0_0_io_A_out_exponent; // @[Array.scala 95:75]
  wire [12:0] array_0_0_io_A_out_fraction; // @[Array.scala 95:75]
  wire  array_0_0_io_B_out_zero; // @[Array.scala 95:75]
  wire  array_0_0_io_B_out_nan; // @[Array.scala 95:75]
  wire  array_0_0_io_B_out_sign; // @[Array.scala 95:75]
  wire [5:0] array_0_0_io_B_out_exponent; // @[Array.scala 95:75]
  wire [12:0] array_0_0_io_B_out_fraction; // @[Array.scala 95:75]
  wire  array_0_0_io_C_out_zero; // @[Array.scala 95:75]
  wire  array_0_0_io_C_out_nan; // @[Array.scala 95:75]
  wire [128:0] array_0_0_io_C_out_number; // @[Array.scala 95:75]
  wire  array_0_0_io_prop_out; // @[Array.scala 95:75]
  wire  array_0_1_clock; // @[Array.scala 95:75]
  wire  array_0_1_io_A_in_zero; // @[Array.scala 95:75]
  wire  array_0_1_io_A_in_nan; // @[Array.scala 95:75]
  wire  array_0_1_io_A_in_sign; // @[Array.scala 95:75]
  wire [5:0] array_0_1_io_A_in_exponent; // @[Array.scala 95:75]
  wire [12:0] array_0_1_io_A_in_fraction; // @[Array.scala 95:75]
  wire  array_0_1_io_B_in_zero; // @[Array.scala 95:75]
  wire  array_0_1_io_B_in_nan; // @[Array.scala 95:75]
  wire  array_0_1_io_B_in_sign; // @[Array.scala 95:75]
  wire [5:0] array_0_1_io_B_in_exponent; // @[Array.scala 95:75]
  wire [12:0] array_0_1_io_B_in_fraction; // @[Array.scala 95:75]
  wire  array_0_1_io_C_in_zero; // @[Array.scala 95:75]
  wire  array_0_1_io_C_in_nan; // @[Array.scala 95:75]
  wire [128:0] array_0_1_io_C_in_number; // @[Array.scala 95:75]
  wire  array_0_1_io_prop_in; // @[Array.scala 95:75]
  wire  array_0_1_io_A_out_zero; // @[Array.scala 95:75]
  wire  array_0_1_io_A_out_nan; // @[Array.scala 95:75]
  wire  array_0_1_io_A_out_sign; // @[Array.scala 95:75]
  wire [5:0] array_0_1_io_A_out_exponent; // @[Array.scala 95:75]
  wire [12:0] array_0_1_io_A_out_fraction; // @[Array.scala 95:75]
  wire  array_0_1_io_B_out_zero; // @[Array.scala 95:75]
  wire  array_0_1_io_B_out_nan; // @[Array.scala 95:75]
  wire  array_0_1_io_B_out_sign; // @[Array.scala 95:75]
  wire [5:0] array_0_1_io_B_out_exponent; // @[Array.scala 95:75]
  wire [12:0] array_0_1_io_B_out_fraction; // @[Array.scala 95:75]
  wire  array_0_1_io_C_out_zero; // @[Array.scala 95:75]
  wire  array_0_1_io_C_out_nan; // @[Array.scala 95:75]
  wire [128:0] array_0_1_io_C_out_number; // @[Array.scala 95:75]
  wire  array_0_1_io_prop_out; // @[Array.scala 95:75]
  wire  array_0_2_clock; // @[Array.scala 95:75]
  wire  array_0_2_io_A_in_zero; // @[Array.scala 95:75]
  wire  array_0_2_io_A_in_nan; // @[Array.scala 95:75]
  wire  array_0_2_io_A_in_sign; // @[Array.scala 95:75]
  wire [5:0] array_0_2_io_A_in_exponent; // @[Array.scala 95:75]
  wire [12:0] array_0_2_io_A_in_fraction; // @[Array.scala 95:75]
  wire  array_0_2_io_B_in_zero; // @[Array.scala 95:75]
  wire  array_0_2_io_B_in_nan; // @[Array.scala 95:75]
  wire  array_0_2_io_B_in_sign; // @[Array.scala 95:75]
  wire [5:0] array_0_2_io_B_in_exponent; // @[Array.scala 95:75]
  wire [12:0] array_0_2_io_B_in_fraction; // @[Array.scala 95:75]
  wire  array_0_2_io_C_in_zero; // @[Array.scala 95:75]
  wire  array_0_2_io_C_in_nan; // @[Array.scala 95:75]
  wire [128:0] array_0_2_io_C_in_number; // @[Array.scala 95:75]
  wire  array_0_2_io_prop_in; // @[Array.scala 95:75]
  wire  array_0_2_io_A_out_zero; // @[Array.scala 95:75]
  wire  array_0_2_io_A_out_nan; // @[Array.scala 95:75]
  wire  array_0_2_io_A_out_sign; // @[Array.scala 95:75]
  wire [5:0] array_0_2_io_A_out_exponent; // @[Array.scala 95:75]
  wire [12:0] array_0_2_io_A_out_fraction; // @[Array.scala 95:75]
  wire  array_0_2_io_B_out_zero; // @[Array.scala 95:75]
  wire  array_0_2_io_B_out_nan; // @[Array.scala 95:75]
  wire  array_0_2_io_B_out_sign; // @[Array.scala 95:75]
  wire [5:0] array_0_2_io_B_out_exponent; // @[Array.scala 95:75]
  wire [12:0] array_0_2_io_B_out_fraction; // @[Array.scala 95:75]
  wire  array_0_2_io_C_out_zero; // @[Array.scala 95:75]
  wire  array_0_2_io_C_out_nan; // @[Array.scala 95:75]
  wire [128:0] array_0_2_io_C_out_number; // @[Array.scala 95:75]
  wire  array_0_2_io_prop_out; // @[Array.scala 95:75]
  wire  array_0_3_clock; // @[Array.scala 95:75]
  wire  array_0_3_io_A_in_zero; // @[Array.scala 95:75]
  wire  array_0_3_io_A_in_nan; // @[Array.scala 95:75]
  wire  array_0_3_io_A_in_sign; // @[Array.scala 95:75]
  wire [5:0] array_0_3_io_A_in_exponent; // @[Array.scala 95:75]
  wire [12:0] array_0_3_io_A_in_fraction; // @[Array.scala 95:75]
  wire  array_0_3_io_B_in_zero; // @[Array.scala 95:75]
  wire  array_0_3_io_B_in_nan; // @[Array.scala 95:75]
  wire  array_0_3_io_B_in_sign; // @[Array.scala 95:75]
  wire [5:0] array_0_3_io_B_in_exponent; // @[Array.scala 95:75]
  wire [12:0] array_0_3_io_B_in_fraction; // @[Array.scala 95:75]
  wire  array_0_3_io_C_in_zero; // @[Array.scala 95:75]
  wire  array_0_3_io_C_in_nan; // @[Array.scala 95:75]
  wire [128:0] array_0_3_io_C_in_number; // @[Array.scala 95:75]
  wire  array_0_3_io_prop_in; // @[Array.scala 95:75]
  wire  array_0_3_io_A_out_zero; // @[Array.scala 95:75]
  wire  array_0_3_io_A_out_nan; // @[Array.scala 95:75]
  wire  array_0_3_io_A_out_sign; // @[Array.scala 95:75]
  wire [5:0] array_0_3_io_A_out_exponent; // @[Array.scala 95:75]
  wire [12:0] array_0_3_io_A_out_fraction; // @[Array.scala 95:75]
  wire  array_0_3_io_B_out_zero; // @[Array.scala 95:75]
  wire  array_0_3_io_B_out_nan; // @[Array.scala 95:75]
  wire  array_0_3_io_B_out_sign; // @[Array.scala 95:75]
  wire [5:0] array_0_3_io_B_out_exponent; // @[Array.scala 95:75]
  wire [12:0] array_0_3_io_B_out_fraction; // @[Array.scala 95:75]
  wire  array_0_3_io_C_out_zero; // @[Array.scala 95:75]
  wire  array_0_3_io_C_out_nan; // @[Array.scala 95:75]
  wire [128:0] array_0_3_io_C_out_number; // @[Array.scala 95:75]
  wire  array_0_3_io_prop_out; // @[Array.scala 95:75]
  wire  array_1_0_clock; // @[Array.scala 95:75]
  wire  array_1_0_io_A_in_zero; // @[Array.scala 95:75]
  wire  array_1_0_io_A_in_nan; // @[Array.scala 95:75]
  wire  array_1_0_io_A_in_sign; // @[Array.scala 95:75]
  wire [5:0] array_1_0_io_A_in_exponent; // @[Array.scala 95:75]
  wire [12:0] array_1_0_io_A_in_fraction; // @[Array.scala 95:75]
  wire  array_1_0_io_B_in_zero; // @[Array.scala 95:75]
  wire  array_1_0_io_B_in_nan; // @[Array.scala 95:75]
  wire  array_1_0_io_B_in_sign; // @[Array.scala 95:75]
  wire [5:0] array_1_0_io_B_in_exponent; // @[Array.scala 95:75]
  wire [12:0] array_1_0_io_B_in_fraction; // @[Array.scala 95:75]
  wire  array_1_0_io_C_in_zero; // @[Array.scala 95:75]
  wire  array_1_0_io_C_in_nan; // @[Array.scala 95:75]
  wire [128:0] array_1_0_io_C_in_number; // @[Array.scala 95:75]
  wire  array_1_0_io_prop_in; // @[Array.scala 95:75]
  wire  array_1_0_io_A_out_zero; // @[Array.scala 95:75]
  wire  array_1_0_io_A_out_nan; // @[Array.scala 95:75]
  wire  array_1_0_io_A_out_sign; // @[Array.scala 95:75]
  wire [5:0] array_1_0_io_A_out_exponent; // @[Array.scala 95:75]
  wire [12:0] array_1_0_io_A_out_fraction; // @[Array.scala 95:75]
  wire  array_1_0_io_B_out_zero; // @[Array.scala 95:75]
  wire  array_1_0_io_B_out_nan; // @[Array.scala 95:75]
  wire  array_1_0_io_B_out_sign; // @[Array.scala 95:75]
  wire [5:0] array_1_0_io_B_out_exponent; // @[Array.scala 95:75]
  wire [12:0] array_1_0_io_B_out_fraction; // @[Array.scala 95:75]
  wire  array_1_0_io_C_out_zero; // @[Array.scala 95:75]
  wire  array_1_0_io_C_out_nan; // @[Array.scala 95:75]
  wire [128:0] array_1_0_io_C_out_number; // @[Array.scala 95:75]
  wire  array_1_0_io_prop_out; // @[Array.scala 95:75]
  wire  array_1_1_clock; // @[Array.scala 95:75]
  wire  array_1_1_io_A_in_zero; // @[Array.scala 95:75]
  wire  array_1_1_io_A_in_nan; // @[Array.scala 95:75]
  wire  array_1_1_io_A_in_sign; // @[Array.scala 95:75]
  wire [5:0] array_1_1_io_A_in_exponent; // @[Array.scala 95:75]
  wire [12:0] array_1_1_io_A_in_fraction; // @[Array.scala 95:75]
  wire  array_1_1_io_B_in_zero; // @[Array.scala 95:75]
  wire  array_1_1_io_B_in_nan; // @[Array.scala 95:75]
  wire  array_1_1_io_B_in_sign; // @[Array.scala 95:75]
  wire [5:0] array_1_1_io_B_in_exponent; // @[Array.scala 95:75]
  wire [12:0] array_1_1_io_B_in_fraction; // @[Array.scala 95:75]
  wire  array_1_1_io_C_in_zero; // @[Array.scala 95:75]
  wire  array_1_1_io_C_in_nan; // @[Array.scala 95:75]
  wire [128:0] array_1_1_io_C_in_number; // @[Array.scala 95:75]
  wire  array_1_1_io_prop_in; // @[Array.scala 95:75]
  wire  array_1_1_io_A_out_zero; // @[Array.scala 95:75]
  wire  array_1_1_io_A_out_nan; // @[Array.scala 95:75]
  wire  array_1_1_io_A_out_sign; // @[Array.scala 95:75]
  wire [5:0] array_1_1_io_A_out_exponent; // @[Array.scala 95:75]
  wire [12:0] array_1_1_io_A_out_fraction; // @[Array.scala 95:75]
  wire  array_1_1_io_B_out_zero; // @[Array.scala 95:75]
  wire  array_1_1_io_B_out_nan; // @[Array.scala 95:75]
  wire  array_1_1_io_B_out_sign; // @[Array.scala 95:75]
  wire [5:0] array_1_1_io_B_out_exponent; // @[Array.scala 95:75]
  wire [12:0] array_1_1_io_B_out_fraction; // @[Array.scala 95:75]
  wire  array_1_1_io_C_out_zero; // @[Array.scala 95:75]
  wire  array_1_1_io_C_out_nan; // @[Array.scala 95:75]
  wire [128:0] array_1_1_io_C_out_number; // @[Array.scala 95:75]
  wire  array_1_1_io_prop_out; // @[Array.scala 95:75]
  wire  array_1_2_clock; // @[Array.scala 95:75]
  wire  array_1_2_io_A_in_zero; // @[Array.scala 95:75]
  wire  array_1_2_io_A_in_nan; // @[Array.scala 95:75]
  wire  array_1_2_io_A_in_sign; // @[Array.scala 95:75]
  wire [5:0] array_1_2_io_A_in_exponent; // @[Array.scala 95:75]
  wire [12:0] array_1_2_io_A_in_fraction; // @[Array.scala 95:75]
  wire  array_1_2_io_B_in_zero; // @[Array.scala 95:75]
  wire  array_1_2_io_B_in_nan; // @[Array.scala 95:75]
  wire  array_1_2_io_B_in_sign; // @[Array.scala 95:75]
  wire [5:0] array_1_2_io_B_in_exponent; // @[Array.scala 95:75]
  wire [12:0] array_1_2_io_B_in_fraction; // @[Array.scala 95:75]
  wire  array_1_2_io_C_in_zero; // @[Array.scala 95:75]
  wire  array_1_2_io_C_in_nan; // @[Array.scala 95:75]
  wire [128:0] array_1_2_io_C_in_number; // @[Array.scala 95:75]
  wire  array_1_2_io_prop_in; // @[Array.scala 95:75]
  wire  array_1_2_io_A_out_zero; // @[Array.scala 95:75]
  wire  array_1_2_io_A_out_nan; // @[Array.scala 95:75]
  wire  array_1_2_io_A_out_sign; // @[Array.scala 95:75]
  wire [5:0] array_1_2_io_A_out_exponent; // @[Array.scala 95:75]
  wire [12:0] array_1_2_io_A_out_fraction; // @[Array.scala 95:75]
  wire  array_1_2_io_B_out_zero; // @[Array.scala 95:75]
  wire  array_1_2_io_B_out_nan; // @[Array.scala 95:75]
  wire  array_1_2_io_B_out_sign; // @[Array.scala 95:75]
  wire [5:0] array_1_2_io_B_out_exponent; // @[Array.scala 95:75]
  wire [12:0] array_1_2_io_B_out_fraction; // @[Array.scala 95:75]
  wire  array_1_2_io_C_out_zero; // @[Array.scala 95:75]
  wire  array_1_2_io_C_out_nan; // @[Array.scala 95:75]
  wire [128:0] array_1_2_io_C_out_number; // @[Array.scala 95:75]
  wire  array_1_2_io_prop_out; // @[Array.scala 95:75]
  wire  array_1_3_clock; // @[Array.scala 95:75]
  wire  array_1_3_io_A_in_zero; // @[Array.scala 95:75]
  wire  array_1_3_io_A_in_nan; // @[Array.scala 95:75]
  wire  array_1_3_io_A_in_sign; // @[Array.scala 95:75]
  wire [5:0] array_1_3_io_A_in_exponent; // @[Array.scala 95:75]
  wire [12:0] array_1_3_io_A_in_fraction; // @[Array.scala 95:75]
  wire  array_1_3_io_B_in_zero; // @[Array.scala 95:75]
  wire  array_1_3_io_B_in_nan; // @[Array.scala 95:75]
  wire  array_1_3_io_B_in_sign; // @[Array.scala 95:75]
  wire [5:0] array_1_3_io_B_in_exponent; // @[Array.scala 95:75]
  wire [12:0] array_1_3_io_B_in_fraction; // @[Array.scala 95:75]
  wire  array_1_3_io_C_in_zero; // @[Array.scala 95:75]
  wire  array_1_3_io_C_in_nan; // @[Array.scala 95:75]
  wire [128:0] array_1_3_io_C_in_number; // @[Array.scala 95:75]
  wire  array_1_3_io_prop_in; // @[Array.scala 95:75]
  wire  array_1_3_io_A_out_zero; // @[Array.scala 95:75]
  wire  array_1_3_io_A_out_nan; // @[Array.scala 95:75]
  wire  array_1_3_io_A_out_sign; // @[Array.scala 95:75]
  wire [5:0] array_1_3_io_A_out_exponent; // @[Array.scala 95:75]
  wire [12:0] array_1_3_io_A_out_fraction; // @[Array.scala 95:75]
  wire  array_1_3_io_B_out_zero; // @[Array.scala 95:75]
  wire  array_1_3_io_B_out_nan; // @[Array.scala 95:75]
  wire  array_1_3_io_B_out_sign; // @[Array.scala 95:75]
  wire [5:0] array_1_3_io_B_out_exponent; // @[Array.scala 95:75]
  wire [12:0] array_1_3_io_B_out_fraction; // @[Array.scala 95:75]
  wire  array_1_3_io_C_out_zero; // @[Array.scala 95:75]
  wire  array_1_3_io_C_out_nan; // @[Array.scala 95:75]
  wire [128:0] array_1_3_io_C_out_number; // @[Array.scala 95:75]
  wire  array_1_3_io_prop_out; // @[Array.scala 95:75]
  wire  array_2_0_clock; // @[Array.scala 95:75]
  wire  array_2_0_io_A_in_zero; // @[Array.scala 95:75]
  wire  array_2_0_io_A_in_nan; // @[Array.scala 95:75]
  wire  array_2_0_io_A_in_sign; // @[Array.scala 95:75]
  wire [5:0] array_2_0_io_A_in_exponent; // @[Array.scala 95:75]
  wire [12:0] array_2_0_io_A_in_fraction; // @[Array.scala 95:75]
  wire  array_2_0_io_B_in_zero; // @[Array.scala 95:75]
  wire  array_2_0_io_B_in_nan; // @[Array.scala 95:75]
  wire  array_2_0_io_B_in_sign; // @[Array.scala 95:75]
  wire [5:0] array_2_0_io_B_in_exponent; // @[Array.scala 95:75]
  wire [12:0] array_2_0_io_B_in_fraction; // @[Array.scala 95:75]
  wire  array_2_0_io_C_in_zero; // @[Array.scala 95:75]
  wire  array_2_0_io_C_in_nan; // @[Array.scala 95:75]
  wire [128:0] array_2_0_io_C_in_number; // @[Array.scala 95:75]
  wire  array_2_0_io_prop_in; // @[Array.scala 95:75]
  wire  array_2_0_io_A_out_zero; // @[Array.scala 95:75]
  wire  array_2_0_io_A_out_nan; // @[Array.scala 95:75]
  wire  array_2_0_io_A_out_sign; // @[Array.scala 95:75]
  wire [5:0] array_2_0_io_A_out_exponent; // @[Array.scala 95:75]
  wire [12:0] array_2_0_io_A_out_fraction; // @[Array.scala 95:75]
  wire  array_2_0_io_B_out_zero; // @[Array.scala 95:75]
  wire  array_2_0_io_B_out_nan; // @[Array.scala 95:75]
  wire  array_2_0_io_B_out_sign; // @[Array.scala 95:75]
  wire [5:0] array_2_0_io_B_out_exponent; // @[Array.scala 95:75]
  wire [12:0] array_2_0_io_B_out_fraction; // @[Array.scala 95:75]
  wire  array_2_0_io_C_out_zero; // @[Array.scala 95:75]
  wire  array_2_0_io_C_out_nan; // @[Array.scala 95:75]
  wire [128:0] array_2_0_io_C_out_number; // @[Array.scala 95:75]
  wire  array_2_0_io_prop_out; // @[Array.scala 95:75]
  wire  array_2_1_clock; // @[Array.scala 95:75]
  wire  array_2_1_io_A_in_zero; // @[Array.scala 95:75]
  wire  array_2_1_io_A_in_nan; // @[Array.scala 95:75]
  wire  array_2_1_io_A_in_sign; // @[Array.scala 95:75]
  wire [5:0] array_2_1_io_A_in_exponent; // @[Array.scala 95:75]
  wire [12:0] array_2_1_io_A_in_fraction; // @[Array.scala 95:75]
  wire  array_2_1_io_B_in_zero; // @[Array.scala 95:75]
  wire  array_2_1_io_B_in_nan; // @[Array.scala 95:75]
  wire  array_2_1_io_B_in_sign; // @[Array.scala 95:75]
  wire [5:0] array_2_1_io_B_in_exponent; // @[Array.scala 95:75]
  wire [12:0] array_2_1_io_B_in_fraction; // @[Array.scala 95:75]
  wire  array_2_1_io_C_in_zero; // @[Array.scala 95:75]
  wire  array_2_1_io_C_in_nan; // @[Array.scala 95:75]
  wire [128:0] array_2_1_io_C_in_number; // @[Array.scala 95:75]
  wire  array_2_1_io_prop_in; // @[Array.scala 95:75]
  wire  array_2_1_io_A_out_zero; // @[Array.scala 95:75]
  wire  array_2_1_io_A_out_nan; // @[Array.scala 95:75]
  wire  array_2_1_io_A_out_sign; // @[Array.scala 95:75]
  wire [5:0] array_2_1_io_A_out_exponent; // @[Array.scala 95:75]
  wire [12:0] array_2_1_io_A_out_fraction; // @[Array.scala 95:75]
  wire  array_2_1_io_B_out_zero; // @[Array.scala 95:75]
  wire  array_2_1_io_B_out_nan; // @[Array.scala 95:75]
  wire  array_2_1_io_B_out_sign; // @[Array.scala 95:75]
  wire [5:0] array_2_1_io_B_out_exponent; // @[Array.scala 95:75]
  wire [12:0] array_2_1_io_B_out_fraction; // @[Array.scala 95:75]
  wire  array_2_1_io_C_out_zero; // @[Array.scala 95:75]
  wire  array_2_1_io_C_out_nan; // @[Array.scala 95:75]
  wire [128:0] array_2_1_io_C_out_number; // @[Array.scala 95:75]
  wire  array_2_1_io_prop_out; // @[Array.scala 95:75]
  wire  array_2_2_clock; // @[Array.scala 95:75]
  wire  array_2_2_io_A_in_zero; // @[Array.scala 95:75]
  wire  array_2_2_io_A_in_nan; // @[Array.scala 95:75]
  wire  array_2_2_io_A_in_sign; // @[Array.scala 95:75]
  wire [5:0] array_2_2_io_A_in_exponent; // @[Array.scala 95:75]
  wire [12:0] array_2_2_io_A_in_fraction; // @[Array.scala 95:75]
  wire  array_2_2_io_B_in_zero; // @[Array.scala 95:75]
  wire  array_2_2_io_B_in_nan; // @[Array.scala 95:75]
  wire  array_2_2_io_B_in_sign; // @[Array.scala 95:75]
  wire [5:0] array_2_2_io_B_in_exponent; // @[Array.scala 95:75]
  wire [12:0] array_2_2_io_B_in_fraction; // @[Array.scala 95:75]
  wire  array_2_2_io_C_in_zero; // @[Array.scala 95:75]
  wire  array_2_2_io_C_in_nan; // @[Array.scala 95:75]
  wire [128:0] array_2_2_io_C_in_number; // @[Array.scala 95:75]
  wire  array_2_2_io_prop_in; // @[Array.scala 95:75]
  wire  array_2_2_io_A_out_zero; // @[Array.scala 95:75]
  wire  array_2_2_io_A_out_nan; // @[Array.scala 95:75]
  wire  array_2_2_io_A_out_sign; // @[Array.scala 95:75]
  wire [5:0] array_2_2_io_A_out_exponent; // @[Array.scala 95:75]
  wire [12:0] array_2_2_io_A_out_fraction; // @[Array.scala 95:75]
  wire  array_2_2_io_B_out_zero; // @[Array.scala 95:75]
  wire  array_2_2_io_B_out_nan; // @[Array.scala 95:75]
  wire  array_2_2_io_B_out_sign; // @[Array.scala 95:75]
  wire [5:0] array_2_2_io_B_out_exponent; // @[Array.scala 95:75]
  wire [12:0] array_2_2_io_B_out_fraction; // @[Array.scala 95:75]
  wire  array_2_2_io_C_out_zero; // @[Array.scala 95:75]
  wire  array_2_2_io_C_out_nan; // @[Array.scala 95:75]
  wire [128:0] array_2_2_io_C_out_number; // @[Array.scala 95:75]
  wire  array_2_2_io_prop_out; // @[Array.scala 95:75]
  wire  array_2_3_clock; // @[Array.scala 95:75]
  wire  array_2_3_io_A_in_zero; // @[Array.scala 95:75]
  wire  array_2_3_io_A_in_nan; // @[Array.scala 95:75]
  wire  array_2_3_io_A_in_sign; // @[Array.scala 95:75]
  wire [5:0] array_2_3_io_A_in_exponent; // @[Array.scala 95:75]
  wire [12:0] array_2_3_io_A_in_fraction; // @[Array.scala 95:75]
  wire  array_2_3_io_B_in_zero; // @[Array.scala 95:75]
  wire  array_2_3_io_B_in_nan; // @[Array.scala 95:75]
  wire  array_2_3_io_B_in_sign; // @[Array.scala 95:75]
  wire [5:0] array_2_3_io_B_in_exponent; // @[Array.scala 95:75]
  wire [12:0] array_2_3_io_B_in_fraction; // @[Array.scala 95:75]
  wire  array_2_3_io_C_in_zero; // @[Array.scala 95:75]
  wire  array_2_3_io_C_in_nan; // @[Array.scala 95:75]
  wire [128:0] array_2_3_io_C_in_number; // @[Array.scala 95:75]
  wire  array_2_3_io_prop_in; // @[Array.scala 95:75]
  wire  array_2_3_io_A_out_zero; // @[Array.scala 95:75]
  wire  array_2_3_io_A_out_nan; // @[Array.scala 95:75]
  wire  array_2_3_io_A_out_sign; // @[Array.scala 95:75]
  wire [5:0] array_2_3_io_A_out_exponent; // @[Array.scala 95:75]
  wire [12:0] array_2_3_io_A_out_fraction; // @[Array.scala 95:75]
  wire  array_2_3_io_B_out_zero; // @[Array.scala 95:75]
  wire  array_2_3_io_B_out_nan; // @[Array.scala 95:75]
  wire  array_2_3_io_B_out_sign; // @[Array.scala 95:75]
  wire [5:0] array_2_3_io_B_out_exponent; // @[Array.scala 95:75]
  wire [12:0] array_2_3_io_B_out_fraction; // @[Array.scala 95:75]
  wire  array_2_3_io_C_out_zero; // @[Array.scala 95:75]
  wire  array_2_3_io_C_out_nan; // @[Array.scala 95:75]
  wire [128:0] array_2_3_io_C_out_number; // @[Array.scala 95:75]
  wire  array_2_3_io_prop_out; // @[Array.scala 95:75]
  wire  array_3_0_clock; // @[Array.scala 95:75]
  wire  array_3_0_io_A_in_zero; // @[Array.scala 95:75]
  wire  array_3_0_io_A_in_nan; // @[Array.scala 95:75]
  wire  array_3_0_io_A_in_sign; // @[Array.scala 95:75]
  wire [5:0] array_3_0_io_A_in_exponent; // @[Array.scala 95:75]
  wire [12:0] array_3_0_io_A_in_fraction; // @[Array.scala 95:75]
  wire  array_3_0_io_B_in_zero; // @[Array.scala 95:75]
  wire  array_3_0_io_B_in_nan; // @[Array.scala 95:75]
  wire  array_3_0_io_B_in_sign; // @[Array.scala 95:75]
  wire [5:0] array_3_0_io_B_in_exponent; // @[Array.scala 95:75]
  wire [12:0] array_3_0_io_B_in_fraction; // @[Array.scala 95:75]
  wire  array_3_0_io_C_in_zero; // @[Array.scala 95:75]
  wire  array_3_0_io_C_in_nan; // @[Array.scala 95:75]
  wire [128:0] array_3_0_io_C_in_number; // @[Array.scala 95:75]
  wire  array_3_0_io_prop_in; // @[Array.scala 95:75]
  wire  array_3_0_io_A_out_zero; // @[Array.scala 95:75]
  wire  array_3_0_io_A_out_nan; // @[Array.scala 95:75]
  wire  array_3_0_io_A_out_sign; // @[Array.scala 95:75]
  wire [5:0] array_3_0_io_A_out_exponent; // @[Array.scala 95:75]
  wire [12:0] array_3_0_io_A_out_fraction; // @[Array.scala 95:75]
  wire  array_3_0_io_B_out_zero; // @[Array.scala 95:75]
  wire  array_3_0_io_B_out_nan; // @[Array.scala 95:75]
  wire  array_3_0_io_B_out_sign; // @[Array.scala 95:75]
  wire [5:0] array_3_0_io_B_out_exponent; // @[Array.scala 95:75]
  wire [12:0] array_3_0_io_B_out_fraction; // @[Array.scala 95:75]
  wire  array_3_0_io_C_out_zero; // @[Array.scala 95:75]
  wire  array_3_0_io_C_out_nan; // @[Array.scala 95:75]
  wire [128:0] array_3_0_io_C_out_number; // @[Array.scala 95:75]
  wire  array_3_0_io_prop_out; // @[Array.scala 95:75]
  wire  array_3_1_clock; // @[Array.scala 95:75]
  wire  array_3_1_io_A_in_zero; // @[Array.scala 95:75]
  wire  array_3_1_io_A_in_nan; // @[Array.scala 95:75]
  wire  array_3_1_io_A_in_sign; // @[Array.scala 95:75]
  wire [5:0] array_3_1_io_A_in_exponent; // @[Array.scala 95:75]
  wire [12:0] array_3_1_io_A_in_fraction; // @[Array.scala 95:75]
  wire  array_3_1_io_B_in_zero; // @[Array.scala 95:75]
  wire  array_3_1_io_B_in_nan; // @[Array.scala 95:75]
  wire  array_3_1_io_B_in_sign; // @[Array.scala 95:75]
  wire [5:0] array_3_1_io_B_in_exponent; // @[Array.scala 95:75]
  wire [12:0] array_3_1_io_B_in_fraction; // @[Array.scala 95:75]
  wire  array_3_1_io_C_in_zero; // @[Array.scala 95:75]
  wire  array_3_1_io_C_in_nan; // @[Array.scala 95:75]
  wire [128:0] array_3_1_io_C_in_number; // @[Array.scala 95:75]
  wire  array_3_1_io_prop_in; // @[Array.scala 95:75]
  wire  array_3_1_io_A_out_zero; // @[Array.scala 95:75]
  wire  array_3_1_io_A_out_nan; // @[Array.scala 95:75]
  wire  array_3_1_io_A_out_sign; // @[Array.scala 95:75]
  wire [5:0] array_3_1_io_A_out_exponent; // @[Array.scala 95:75]
  wire [12:0] array_3_1_io_A_out_fraction; // @[Array.scala 95:75]
  wire  array_3_1_io_B_out_zero; // @[Array.scala 95:75]
  wire  array_3_1_io_B_out_nan; // @[Array.scala 95:75]
  wire  array_3_1_io_B_out_sign; // @[Array.scala 95:75]
  wire [5:0] array_3_1_io_B_out_exponent; // @[Array.scala 95:75]
  wire [12:0] array_3_1_io_B_out_fraction; // @[Array.scala 95:75]
  wire  array_3_1_io_C_out_zero; // @[Array.scala 95:75]
  wire  array_3_1_io_C_out_nan; // @[Array.scala 95:75]
  wire [128:0] array_3_1_io_C_out_number; // @[Array.scala 95:75]
  wire  array_3_1_io_prop_out; // @[Array.scala 95:75]
  wire  array_3_2_clock; // @[Array.scala 95:75]
  wire  array_3_2_io_A_in_zero; // @[Array.scala 95:75]
  wire  array_3_2_io_A_in_nan; // @[Array.scala 95:75]
  wire  array_3_2_io_A_in_sign; // @[Array.scala 95:75]
  wire [5:0] array_3_2_io_A_in_exponent; // @[Array.scala 95:75]
  wire [12:0] array_3_2_io_A_in_fraction; // @[Array.scala 95:75]
  wire  array_3_2_io_B_in_zero; // @[Array.scala 95:75]
  wire  array_3_2_io_B_in_nan; // @[Array.scala 95:75]
  wire  array_3_2_io_B_in_sign; // @[Array.scala 95:75]
  wire [5:0] array_3_2_io_B_in_exponent; // @[Array.scala 95:75]
  wire [12:0] array_3_2_io_B_in_fraction; // @[Array.scala 95:75]
  wire  array_3_2_io_C_in_zero; // @[Array.scala 95:75]
  wire  array_3_2_io_C_in_nan; // @[Array.scala 95:75]
  wire [128:0] array_3_2_io_C_in_number; // @[Array.scala 95:75]
  wire  array_3_2_io_prop_in; // @[Array.scala 95:75]
  wire  array_3_2_io_A_out_zero; // @[Array.scala 95:75]
  wire  array_3_2_io_A_out_nan; // @[Array.scala 95:75]
  wire  array_3_2_io_A_out_sign; // @[Array.scala 95:75]
  wire [5:0] array_3_2_io_A_out_exponent; // @[Array.scala 95:75]
  wire [12:0] array_3_2_io_A_out_fraction; // @[Array.scala 95:75]
  wire  array_3_2_io_B_out_zero; // @[Array.scala 95:75]
  wire  array_3_2_io_B_out_nan; // @[Array.scala 95:75]
  wire  array_3_2_io_B_out_sign; // @[Array.scala 95:75]
  wire [5:0] array_3_2_io_B_out_exponent; // @[Array.scala 95:75]
  wire [12:0] array_3_2_io_B_out_fraction; // @[Array.scala 95:75]
  wire  array_3_2_io_C_out_zero; // @[Array.scala 95:75]
  wire  array_3_2_io_C_out_nan; // @[Array.scala 95:75]
  wire [128:0] array_3_2_io_C_out_number; // @[Array.scala 95:75]
  wire  array_3_2_io_prop_out; // @[Array.scala 95:75]
  wire  array_3_3_clock; // @[Array.scala 95:75]
  wire  array_3_3_io_A_in_zero; // @[Array.scala 95:75]
  wire  array_3_3_io_A_in_nan; // @[Array.scala 95:75]
  wire  array_3_3_io_A_in_sign; // @[Array.scala 95:75]
  wire [5:0] array_3_3_io_A_in_exponent; // @[Array.scala 95:75]
  wire [12:0] array_3_3_io_A_in_fraction; // @[Array.scala 95:75]
  wire  array_3_3_io_B_in_zero; // @[Array.scala 95:75]
  wire  array_3_3_io_B_in_nan; // @[Array.scala 95:75]
  wire  array_3_3_io_B_in_sign; // @[Array.scala 95:75]
  wire [5:0] array_3_3_io_B_in_exponent; // @[Array.scala 95:75]
  wire [12:0] array_3_3_io_B_in_fraction; // @[Array.scala 95:75]
  wire  array_3_3_io_C_in_zero; // @[Array.scala 95:75]
  wire  array_3_3_io_C_in_nan; // @[Array.scala 95:75]
  wire [128:0] array_3_3_io_C_in_number; // @[Array.scala 95:75]
  wire  array_3_3_io_prop_in; // @[Array.scala 95:75]
  wire  array_3_3_io_A_out_zero; // @[Array.scala 95:75]
  wire  array_3_3_io_A_out_nan; // @[Array.scala 95:75]
  wire  array_3_3_io_A_out_sign; // @[Array.scala 95:75]
  wire [5:0] array_3_3_io_A_out_exponent; // @[Array.scala 95:75]
  wire [12:0] array_3_3_io_A_out_fraction; // @[Array.scala 95:75]
  wire  array_3_3_io_B_out_zero; // @[Array.scala 95:75]
  wire  array_3_3_io_B_out_nan; // @[Array.scala 95:75]
  wire  array_3_3_io_B_out_sign; // @[Array.scala 95:75]
  wire [5:0] array_3_3_io_B_out_exponent; // @[Array.scala 95:75]
  wire [12:0] array_3_3_io_B_out_fraction; // @[Array.scala 95:75]
  wire  array_3_3_io_C_out_zero; // @[Array.scala 95:75]
  wire  array_3_3_io_C_out_nan; // @[Array.scala 95:75]
  wire [128:0] array_3_3_io_C_out_number; // @[Array.scala 95:75]
  wire  array_3_3_io_prop_out; // @[Array.scala 95:75]
  wire [15:0] A_convert_0_io_in; // @[Array.scala 98:76]
  wire  A_convert_0_io_out_zero; // @[Array.scala 98:76]
  wire  A_convert_0_io_out_nan; // @[Array.scala 98:76]
  wire  A_convert_0_io_out_sign; // @[Array.scala 98:76]
  wire [5:0] A_convert_0_io_out_exponent; // @[Array.scala 98:76]
  wire [12:0] A_convert_0_io_out_fraction; // @[Array.scala 98:76]
  wire [15:0] A_convert_1_io_in; // @[Array.scala 98:76]
  wire  A_convert_1_io_out_zero; // @[Array.scala 98:76]
  wire  A_convert_1_io_out_nan; // @[Array.scala 98:76]
  wire  A_convert_1_io_out_sign; // @[Array.scala 98:76]
  wire [5:0] A_convert_1_io_out_exponent; // @[Array.scala 98:76]
  wire [12:0] A_convert_1_io_out_fraction; // @[Array.scala 98:76]
  wire [15:0] A_convert_2_io_in; // @[Array.scala 98:76]
  wire  A_convert_2_io_out_zero; // @[Array.scala 98:76]
  wire  A_convert_2_io_out_nan; // @[Array.scala 98:76]
  wire  A_convert_2_io_out_sign; // @[Array.scala 98:76]
  wire [5:0] A_convert_2_io_out_exponent; // @[Array.scala 98:76]
  wire [12:0] A_convert_2_io_out_fraction; // @[Array.scala 98:76]
  wire [15:0] A_convert_3_io_in; // @[Array.scala 98:76]
  wire  A_convert_3_io_out_zero; // @[Array.scala 98:76]
  wire  A_convert_3_io_out_nan; // @[Array.scala 98:76]
  wire  A_convert_3_io_out_sign; // @[Array.scala 98:76]
  wire [5:0] A_convert_3_io_out_exponent; // @[Array.scala 98:76]
  wire [12:0] A_convert_3_io_out_fraction; // @[Array.scala 98:76]
  wire [15:0] B_convert_0_io_in; // @[Array.scala 99:76]
  wire  B_convert_0_io_out_zero; // @[Array.scala 99:76]
  wire  B_convert_0_io_out_nan; // @[Array.scala 99:76]
  wire  B_convert_0_io_out_sign; // @[Array.scala 99:76]
  wire [5:0] B_convert_0_io_out_exponent; // @[Array.scala 99:76]
  wire [12:0] B_convert_0_io_out_fraction; // @[Array.scala 99:76]
  wire [15:0] B_convert_1_io_in; // @[Array.scala 99:76]
  wire  B_convert_1_io_out_zero; // @[Array.scala 99:76]
  wire  B_convert_1_io_out_nan; // @[Array.scala 99:76]
  wire  B_convert_1_io_out_sign; // @[Array.scala 99:76]
  wire [5:0] B_convert_1_io_out_exponent; // @[Array.scala 99:76]
  wire [12:0] B_convert_1_io_out_fraction; // @[Array.scala 99:76]
  wire [15:0] B_convert_2_io_in; // @[Array.scala 99:76]
  wire  B_convert_2_io_out_zero; // @[Array.scala 99:76]
  wire  B_convert_2_io_out_nan; // @[Array.scala 99:76]
  wire  B_convert_2_io_out_sign; // @[Array.scala 99:76]
  wire [5:0] B_convert_2_io_out_exponent; // @[Array.scala 99:76]
  wire [12:0] B_convert_2_io_out_fraction; // @[Array.scala 99:76]
  wire [15:0] B_convert_3_io_in; // @[Array.scala 99:76]
  wire  B_convert_3_io_out_zero; // @[Array.scala 99:76]
  wire  B_convert_3_io_out_nan; // @[Array.scala 99:76]
  wire  B_convert_3_io_out_sign; // @[Array.scala 99:76]
  wire [5:0] B_convert_3_io_out_exponent; // @[Array.scala 99:76]
  wire [12:0] B_convert_3_io_out_fraction; // @[Array.scala 99:76]
  logTile array_0_0 ( // @[Array.scala 95:75]
    .clock(array_0_0_clock),
    .io_A_in_zero(array_0_0_io_A_in_zero),
    .io_A_in_nan(array_0_0_io_A_in_nan),
    .io_A_in_sign(array_0_0_io_A_in_sign),
    .io_A_in_exponent(array_0_0_io_A_in_exponent),
    .io_A_in_fraction(array_0_0_io_A_in_fraction),
    .io_B_in_zero(array_0_0_io_B_in_zero),
    .io_B_in_nan(array_0_0_io_B_in_nan),
    .io_B_in_sign(array_0_0_io_B_in_sign),
    .io_B_in_exponent(array_0_0_io_B_in_exponent),
    .io_B_in_fraction(array_0_0_io_B_in_fraction),
    .io_C_in_zero(array_0_0_io_C_in_zero),
    .io_C_in_nan(array_0_0_io_C_in_nan),
    .io_C_in_number(array_0_0_io_C_in_number),
    .io_prop_in(array_0_0_io_prop_in),
    .io_A_out_zero(array_0_0_io_A_out_zero),
    .io_A_out_nan(array_0_0_io_A_out_nan),
    .io_A_out_sign(array_0_0_io_A_out_sign),
    .io_A_out_exponent(array_0_0_io_A_out_exponent),
    .io_A_out_fraction(array_0_0_io_A_out_fraction),
    .io_B_out_zero(array_0_0_io_B_out_zero),
    .io_B_out_nan(array_0_0_io_B_out_nan),
    .io_B_out_sign(array_0_0_io_B_out_sign),
    .io_B_out_exponent(array_0_0_io_B_out_exponent),
    .io_B_out_fraction(array_0_0_io_B_out_fraction),
    .io_C_out_zero(array_0_0_io_C_out_zero),
    .io_C_out_nan(array_0_0_io_C_out_nan),
    .io_C_out_number(array_0_0_io_C_out_number),
    .io_prop_out(array_0_0_io_prop_out)
  );
  logTile array_0_1 ( // @[Array.scala 95:75]
    .clock(array_0_1_clock),
    .io_A_in_zero(array_0_1_io_A_in_zero),
    .io_A_in_nan(array_0_1_io_A_in_nan),
    .io_A_in_sign(array_0_1_io_A_in_sign),
    .io_A_in_exponent(array_0_1_io_A_in_exponent),
    .io_A_in_fraction(array_0_1_io_A_in_fraction),
    .io_B_in_zero(array_0_1_io_B_in_zero),
    .io_B_in_nan(array_0_1_io_B_in_nan),
    .io_B_in_sign(array_0_1_io_B_in_sign),
    .io_B_in_exponent(array_0_1_io_B_in_exponent),
    .io_B_in_fraction(array_0_1_io_B_in_fraction),
    .io_C_in_zero(array_0_1_io_C_in_zero),
    .io_C_in_nan(array_0_1_io_C_in_nan),
    .io_C_in_number(array_0_1_io_C_in_number),
    .io_prop_in(array_0_1_io_prop_in),
    .io_A_out_zero(array_0_1_io_A_out_zero),
    .io_A_out_nan(array_0_1_io_A_out_nan),
    .io_A_out_sign(array_0_1_io_A_out_sign),
    .io_A_out_exponent(array_0_1_io_A_out_exponent),
    .io_A_out_fraction(array_0_1_io_A_out_fraction),
    .io_B_out_zero(array_0_1_io_B_out_zero),
    .io_B_out_nan(array_0_1_io_B_out_nan),
    .io_B_out_sign(array_0_1_io_B_out_sign),
    .io_B_out_exponent(array_0_1_io_B_out_exponent),
    .io_B_out_fraction(array_0_1_io_B_out_fraction),
    .io_C_out_zero(array_0_1_io_C_out_zero),
    .io_C_out_nan(array_0_1_io_C_out_nan),
    .io_C_out_number(array_0_1_io_C_out_number),
    .io_prop_out(array_0_1_io_prop_out)
  );
  logTile array_0_2 ( // @[Array.scala 95:75]
    .clock(array_0_2_clock),
    .io_A_in_zero(array_0_2_io_A_in_zero),
    .io_A_in_nan(array_0_2_io_A_in_nan),
    .io_A_in_sign(array_0_2_io_A_in_sign),
    .io_A_in_exponent(array_0_2_io_A_in_exponent),
    .io_A_in_fraction(array_0_2_io_A_in_fraction),
    .io_B_in_zero(array_0_2_io_B_in_zero),
    .io_B_in_nan(array_0_2_io_B_in_nan),
    .io_B_in_sign(array_0_2_io_B_in_sign),
    .io_B_in_exponent(array_0_2_io_B_in_exponent),
    .io_B_in_fraction(array_0_2_io_B_in_fraction),
    .io_C_in_zero(array_0_2_io_C_in_zero),
    .io_C_in_nan(array_0_2_io_C_in_nan),
    .io_C_in_number(array_0_2_io_C_in_number),
    .io_prop_in(array_0_2_io_prop_in),
    .io_A_out_zero(array_0_2_io_A_out_zero),
    .io_A_out_nan(array_0_2_io_A_out_nan),
    .io_A_out_sign(array_0_2_io_A_out_sign),
    .io_A_out_exponent(array_0_2_io_A_out_exponent),
    .io_A_out_fraction(array_0_2_io_A_out_fraction),
    .io_B_out_zero(array_0_2_io_B_out_zero),
    .io_B_out_nan(array_0_2_io_B_out_nan),
    .io_B_out_sign(array_0_2_io_B_out_sign),
    .io_B_out_exponent(array_0_2_io_B_out_exponent),
    .io_B_out_fraction(array_0_2_io_B_out_fraction),
    .io_C_out_zero(array_0_2_io_C_out_zero),
    .io_C_out_nan(array_0_2_io_C_out_nan),
    .io_C_out_number(array_0_2_io_C_out_number),
    .io_prop_out(array_0_2_io_prop_out)
  );
  logTile array_0_3 ( // @[Array.scala 95:75]
    .clock(array_0_3_clock),
    .io_A_in_zero(array_0_3_io_A_in_zero),
    .io_A_in_nan(array_0_3_io_A_in_nan),
    .io_A_in_sign(array_0_3_io_A_in_sign),
    .io_A_in_exponent(array_0_3_io_A_in_exponent),
    .io_A_in_fraction(array_0_3_io_A_in_fraction),
    .io_B_in_zero(array_0_3_io_B_in_zero),
    .io_B_in_nan(array_0_3_io_B_in_nan),
    .io_B_in_sign(array_0_3_io_B_in_sign),
    .io_B_in_exponent(array_0_3_io_B_in_exponent),
    .io_B_in_fraction(array_0_3_io_B_in_fraction),
    .io_C_in_zero(array_0_3_io_C_in_zero),
    .io_C_in_nan(array_0_3_io_C_in_nan),
    .io_C_in_number(array_0_3_io_C_in_number),
    .io_prop_in(array_0_3_io_prop_in),
    .io_A_out_zero(array_0_3_io_A_out_zero),
    .io_A_out_nan(array_0_3_io_A_out_nan),
    .io_A_out_sign(array_0_3_io_A_out_sign),
    .io_A_out_exponent(array_0_3_io_A_out_exponent),
    .io_A_out_fraction(array_0_3_io_A_out_fraction),
    .io_B_out_zero(array_0_3_io_B_out_zero),
    .io_B_out_nan(array_0_3_io_B_out_nan),
    .io_B_out_sign(array_0_3_io_B_out_sign),
    .io_B_out_exponent(array_0_3_io_B_out_exponent),
    .io_B_out_fraction(array_0_3_io_B_out_fraction),
    .io_C_out_zero(array_0_3_io_C_out_zero),
    .io_C_out_nan(array_0_3_io_C_out_nan),
    .io_C_out_number(array_0_3_io_C_out_number),
    .io_prop_out(array_0_3_io_prop_out)
  );
  logTile array_1_0 ( // @[Array.scala 95:75]
    .clock(array_1_0_clock),
    .io_A_in_zero(array_1_0_io_A_in_zero),
    .io_A_in_nan(array_1_0_io_A_in_nan),
    .io_A_in_sign(array_1_0_io_A_in_sign),
    .io_A_in_exponent(array_1_0_io_A_in_exponent),
    .io_A_in_fraction(array_1_0_io_A_in_fraction),
    .io_B_in_zero(array_1_0_io_B_in_zero),
    .io_B_in_nan(array_1_0_io_B_in_nan),
    .io_B_in_sign(array_1_0_io_B_in_sign),
    .io_B_in_exponent(array_1_0_io_B_in_exponent),
    .io_B_in_fraction(array_1_0_io_B_in_fraction),
    .io_C_in_zero(array_1_0_io_C_in_zero),
    .io_C_in_nan(array_1_0_io_C_in_nan),
    .io_C_in_number(array_1_0_io_C_in_number),
    .io_prop_in(array_1_0_io_prop_in),
    .io_A_out_zero(array_1_0_io_A_out_zero),
    .io_A_out_nan(array_1_0_io_A_out_nan),
    .io_A_out_sign(array_1_0_io_A_out_sign),
    .io_A_out_exponent(array_1_0_io_A_out_exponent),
    .io_A_out_fraction(array_1_0_io_A_out_fraction),
    .io_B_out_zero(array_1_0_io_B_out_zero),
    .io_B_out_nan(array_1_0_io_B_out_nan),
    .io_B_out_sign(array_1_0_io_B_out_sign),
    .io_B_out_exponent(array_1_0_io_B_out_exponent),
    .io_B_out_fraction(array_1_0_io_B_out_fraction),
    .io_C_out_zero(array_1_0_io_C_out_zero),
    .io_C_out_nan(array_1_0_io_C_out_nan),
    .io_C_out_number(array_1_0_io_C_out_number),
    .io_prop_out(array_1_0_io_prop_out)
  );
  logTile array_1_1 ( // @[Array.scala 95:75]
    .clock(array_1_1_clock),
    .io_A_in_zero(array_1_1_io_A_in_zero),
    .io_A_in_nan(array_1_1_io_A_in_nan),
    .io_A_in_sign(array_1_1_io_A_in_sign),
    .io_A_in_exponent(array_1_1_io_A_in_exponent),
    .io_A_in_fraction(array_1_1_io_A_in_fraction),
    .io_B_in_zero(array_1_1_io_B_in_zero),
    .io_B_in_nan(array_1_1_io_B_in_nan),
    .io_B_in_sign(array_1_1_io_B_in_sign),
    .io_B_in_exponent(array_1_1_io_B_in_exponent),
    .io_B_in_fraction(array_1_1_io_B_in_fraction),
    .io_C_in_zero(array_1_1_io_C_in_zero),
    .io_C_in_nan(array_1_1_io_C_in_nan),
    .io_C_in_number(array_1_1_io_C_in_number),
    .io_prop_in(array_1_1_io_prop_in),
    .io_A_out_zero(array_1_1_io_A_out_zero),
    .io_A_out_nan(array_1_1_io_A_out_nan),
    .io_A_out_sign(array_1_1_io_A_out_sign),
    .io_A_out_exponent(array_1_1_io_A_out_exponent),
    .io_A_out_fraction(array_1_1_io_A_out_fraction),
    .io_B_out_zero(array_1_1_io_B_out_zero),
    .io_B_out_nan(array_1_1_io_B_out_nan),
    .io_B_out_sign(array_1_1_io_B_out_sign),
    .io_B_out_exponent(array_1_1_io_B_out_exponent),
    .io_B_out_fraction(array_1_1_io_B_out_fraction),
    .io_C_out_zero(array_1_1_io_C_out_zero),
    .io_C_out_nan(array_1_1_io_C_out_nan),
    .io_C_out_number(array_1_1_io_C_out_number),
    .io_prop_out(array_1_1_io_prop_out)
  );
  logTile array_1_2 ( // @[Array.scala 95:75]
    .clock(array_1_2_clock),
    .io_A_in_zero(array_1_2_io_A_in_zero),
    .io_A_in_nan(array_1_2_io_A_in_nan),
    .io_A_in_sign(array_1_2_io_A_in_sign),
    .io_A_in_exponent(array_1_2_io_A_in_exponent),
    .io_A_in_fraction(array_1_2_io_A_in_fraction),
    .io_B_in_zero(array_1_2_io_B_in_zero),
    .io_B_in_nan(array_1_2_io_B_in_nan),
    .io_B_in_sign(array_1_2_io_B_in_sign),
    .io_B_in_exponent(array_1_2_io_B_in_exponent),
    .io_B_in_fraction(array_1_2_io_B_in_fraction),
    .io_C_in_zero(array_1_2_io_C_in_zero),
    .io_C_in_nan(array_1_2_io_C_in_nan),
    .io_C_in_number(array_1_2_io_C_in_number),
    .io_prop_in(array_1_2_io_prop_in),
    .io_A_out_zero(array_1_2_io_A_out_zero),
    .io_A_out_nan(array_1_2_io_A_out_nan),
    .io_A_out_sign(array_1_2_io_A_out_sign),
    .io_A_out_exponent(array_1_2_io_A_out_exponent),
    .io_A_out_fraction(array_1_2_io_A_out_fraction),
    .io_B_out_zero(array_1_2_io_B_out_zero),
    .io_B_out_nan(array_1_2_io_B_out_nan),
    .io_B_out_sign(array_1_2_io_B_out_sign),
    .io_B_out_exponent(array_1_2_io_B_out_exponent),
    .io_B_out_fraction(array_1_2_io_B_out_fraction),
    .io_C_out_zero(array_1_2_io_C_out_zero),
    .io_C_out_nan(array_1_2_io_C_out_nan),
    .io_C_out_number(array_1_2_io_C_out_number),
    .io_prop_out(array_1_2_io_prop_out)
  );
  logTile array_1_3 ( // @[Array.scala 95:75]
    .clock(array_1_3_clock),
    .io_A_in_zero(array_1_3_io_A_in_zero),
    .io_A_in_nan(array_1_3_io_A_in_nan),
    .io_A_in_sign(array_1_3_io_A_in_sign),
    .io_A_in_exponent(array_1_3_io_A_in_exponent),
    .io_A_in_fraction(array_1_3_io_A_in_fraction),
    .io_B_in_zero(array_1_3_io_B_in_zero),
    .io_B_in_nan(array_1_3_io_B_in_nan),
    .io_B_in_sign(array_1_3_io_B_in_sign),
    .io_B_in_exponent(array_1_3_io_B_in_exponent),
    .io_B_in_fraction(array_1_3_io_B_in_fraction),
    .io_C_in_zero(array_1_3_io_C_in_zero),
    .io_C_in_nan(array_1_3_io_C_in_nan),
    .io_C_in_number(array_1_3_io_C_in_number),
    .io_prop_in(array_1_3_io_prop_in),
    .io_A_out_zero(array_1_3_io_A_out_zero),
    .io_A_out_nan(array_1_3_io_A_out_nan),
    .io_A_out_sign(array_1_3_io_A_out_sign),
    .io_A_out_exponent(array_1_3_io_A_out_exponent),
    .io_A_out_fraction(array_1_3_io_A_out_fraction),
    .io_B_out_zero(array_1_3_io_B_out_zero),
    .io_B_out_nan(array_1_3_io_B_out_nan),
    .io_B_out_sign(array_1_3_io_B_out_sign),
    .io_B_out_exponent(array_1_3_io_B_out_exponent),
    .io_B_out_fraction(array_1_3_io_B_out_fraction),
    .io_C_out_zero(array_1_3_io_C_out_zero),
    .io_C_out_nan(array_1_3_io_C_out_nan),
    .io_C_out_number(array_1_3_io_C_out_number),
    .io_prop_out(array_1_3_io_prop_out)
  );
  logTile array_2_0 ( // @[Array.scala 95:75]
    .clock(array_2_0_clock),
    .io_A_in_zero(array_2_0_io_A_in_zero),
    .io_A_in_nan(array_2_0_io_A_in_nan),
    .io_A_in_sign(array_2_0_io_A_in_sign),
    .io_A_in_exponent(array_2_0_io_A_in_exponent),
    .io_A_in_fraction(array_2_0_io_A_in_fraction),
    .io_B_in_zero(array_2_0_io_B_in_zero),
    .io_B_in_nan(array_2_0_io_B_in_nan),
    .io_B_in_sign(array_2_0_io_B_in_sign),
    .io_B_in_exponent(array_2_0_io_B_in_exponent),
    .io_B_in_fraction(array_2_0_io_B_in_fraction),
    .io_C_in_zero(array_2_0_io_C_in_zero),
    .io_C_in_nan(array_2_0_io_C_in_nan),
    .io_C_in_number(array_2_0_io_C_in_number),
    .io_prop_in(array_2_0_io_prop_in),
    .io_A_out_zero(array_2_0_io_A_out_zero),
    .io_A_out_nan(array_2_0_io_A_out_nan),
    .io_A_out_sign(array_2_0_io_A_out_sign),
    .io_A_out_exponent(array_2_0_io_A_out_exponent),
    .io_A_out_fraction(array_2_0_io_A_out_fraction),
    .io_B_out_zero(array_2_0_io_B_out_zero),
    .io_B_out_nan(array_2_0_io_B_out_nan),
    .io_B_out_sign(array_2_0_io_B_out_sign),
    .io_B_out_exponent(array_2_0_io_B_out_exponent),
    .io_B_out_fraction(array_2_0_io_B_out_fraction),
    .io_C_out_zero(array_2_0_io_C_out_zero),
    .io_C_out_nan(array_2_0_io_C_out_nan),
    .io_C_out_number(array_2_0_io_C_out_number),
    .io_prop_out(array_2_0_io_prop_out)
  );
  logTile array_2_1 ( // @[Array.scala 95:75]
    .clock(array_2_1_clock),
    .io_A_in_zero(array_2_1_io_A_in_zero),
    .io_A_in_nan(array_2_1_io_A_in_nan),
    .io_A_in_sign(array_2_1_io_A_in_sign),
    .io_A_in_exponent(array_2_1_io_A_in_exponent),
    .io_A_in_fraction(array_2_1_io_A_in_fraction),
    .io_B_in_zero(array_2_1_io_B_in_zero),
    .io_B_in_nan(array_2_1_io_B_in_nan),
    .io_B_in_sign(array_2_1_io_B_in_sign),
    .io_B_in_exponent(array_2_1_io_B_in_exponent),
    .io_B_in_fraction(array_2_1_io_B_in_fraction),
    .io_C_in_zero(array_2_1_io_C_in_zero),
    .io_C_in_nan(array_2_1_io_C_in_nan),
    .io_C_in_number(array_2_1_io_C_in_number),
    .io_prop_in(array_2_1_io_prop_in),
    .io_A_out_zero(array_2_1_io_A_out_zero),
    .io_A_out_nan(array_2_1_io_A_out_nan),
    .io_A_out_sign(array_2_1_io_A_out_sign),
    .io_A_out_exponent(array_2_1_io_A_out_exponent),
    .io_A_out_fraction(array_2_1_io_A_out_fraction),
    .io_B_out_zero(array_2_1_io_B_out_zero),
    .io_B_out_nan(array_2_1_io_B_out_nan),
    .io_B_out_sign(array_2_1_io_B_out_sign),
    .io_B_out_exponent(array_2_1_io_B_out_exponent),
    .io_B_out_fraction(array_2_1_io_B_out_fraction),
    .io_C_out_zero(array_2_1_io_C_out_zero),
    .io_C_out_nan(array_2_1_io_C_out_nan),
    .io_C_out_number(array_2_1_io_C_out_number),
    .io_prop_out(array_2_1_io_prop_out)
  );
  logTile array_2_2 ( // @[Array.scala 95:75]
    .clock(array_2_2_clock),
    .io_A_in_zero(array_2_2_io_A_in_zero),
    .io_A_in_nan(array_2_2_io_A_in_nan),
    .io_A_in_sign(array_2_2_io_A_in_sign),
    .io_A_in_exponent(array_2_2_io_A_in_exponent),
    .io_A_in_fraction(array_2_2_io_A_in_fraction),
    .io_B_in_zero(array_2_2_io_B_in_zero),
    .io_B_in_nan(array_2_2_io_B_in_nan),
    .io_B_in_sign(array_2_2_io_B_in_sign),
    .io_B_in_exponent(array_2_2_io_B_in_exponent),
    .io_B_in_fraction(array_2_2_io_B_in_fraction),
    .io_C_in_zero(array_2_2_io_C_in_zero),
    .io_C_in_nan(array_2_2_io_C_in_nan),
    .io_C_in_number(array_2_2_io_C_in_number),
    .io_prop_in(array_2_2_io_prop_in),
    .io_A_out_zero(array_2_2_io_A_out_zero),
    .io_A_out_nan(array_2_2_io_A_out_nan),
    .io_A_out_sign(array_2_2_io_A_out_sign),
    .io_A_out_exponent(array_2_2_io_A_out_exponent),
    .io_A_out_fraction(array_2_2_io_A_out_fraction),
    .io_B_out_zero(array_2_2_io_B_out_zero),
    .io_B_out_nan(array_2_2_io_B_out_nan),
    .io_B_out_sign(array_2_2_io_B_out_sign),
    .io_B_out_exponent(array_2_2_io_B_out_exponent),
    .io_B_out_fraction(array_2_2_io_B_out_fraction),
    .io_C_out_zero(array_2_2_io_C_out_zero),
    .io_C_out_nan(array_2_2_io_C_out_nan),
    .io_C_out_number(array_2_2_io_C_out_number),
    .io_prop_out(array_2_2_io_prop_out)
  );
  logTile array_2_3 ( // @[Array.scala 95:75]
    .clock(array_2_3_clock),
    .io_A_in_zero(array_2_3_io_A_in_zero),
    .io_A_in_nan(array_2_3_io_A_in_nan),
    .io_A_in_sign(array_2_3_io_A_in_sign),
    .io_A_in_exponent(array_2_3_io_A_in_exponent),
    .io_A_in_fraction(array_2_3_io_A_in_fraction),
    .io_B_in_zero(array_2_3_io_B_in_zero),
    .io_B_in_nan(array_2_3_io_B_in_nan),
    .io_B_in_sign(array_2_3_io_B_in_sign),
    .io_B_in_exponent(array_2_3_io_B_in_exponent),
    .io_B_in_fraction(array_2_3_io_B_in_fraction),
    .io_C_in_zero(array_2_3_io_C_in_zero),
    .io_C_in_nan(array_2_3_io_C_in_nan),
    .io_C_in_number(array_2_3_io_C_in_number),
    .io_prop_in(array_2_3_io_prop_in),
    .io_A_out_zero(array_2_3_io_A_out_zero),
    .io_A_out_nan(array_2_3_io_A_out_nan),
    .io_A_out_sign(array_2_3_io_A_out_sign),
    .io_A_out_exponent(array_2_3_io_A_out_exponent),
    .io_A_out_fraction(array_2_3_io_A_out_fraction),
    .io_B_out_zero(array_2_3_io_B_out_zero),
    .io_B_out_nan(array_2_3_io_B_out_nan),
    .io_B_out_sign(array_2_3_io_B_out_sign),
    .io_B_out_exponent(array_2_3_io_B_out_exponent),
    .io_B_out_fraction(array_2_3_io_B_out_fraction),
    .io_C_out_zero(array_2_3_io_C_out_zero),
    .io_C_out_nan(array_2_3_io_C_out_nan),
    .io_C_out_number(array_2_3_io_C_out_number),
    .io_prop_out(array_2_3_io_prop_out)
  );
  logTile array_3_0 ( // @[Array.scala 95:75]
    .clock(array_3_0_clock),
    .io_A_in_zero(array_3_0_io_A_in_zero),
    .io_A_in_nan(array_3_0_io_A_in_nan),
    .io_A_in_sign(array_3_0_io_A_in_sign),
    .io_A_in_exponent(array_3_0_io_A_in_exponent),
    .io_A_in_fraction(array_3_0_io_A_in_fraction),
    .io_B_in_zero(array_3_0_io_B_in_zero),
    .io_B_in_nan(array_3_0_io_B_in_nan),
    .io_B_in_sign(array_3_0_io_B_in_sign),
    .io_B_in_exponent(array_3_0_io_B_in_exponent),
    .io_B_in_fraction(array_3_0_io_B_in_fraction),
    .io_C_in_zero(array_3_0_io_C_in_zero),
    .io_C_in_nan(array_3_0_io_C_in_nan),
    .io_C_in_number(array_3_0_io_C_in_number),
    .io_prop_in(array_3_0_io_prop_in),
    .io_A_out_zero(array_3_0_io_A_out_zero),
    .io_A_out_nan(array_3_0_io_A_out_nan),
    .io_A_out_sign(array_3_0_io_A_out_sign),
    .io_A_out_exponent(array_3_0_io_A_out_exponent),
    .io_A_out_fraction(array_3_0_io_A_out_fraction),
    .io_B_out_zero(array_3_0_io_B_out_zero),
    .io_B_out_nan(array_3_0_io_B_out_nan),
    .io_B_out_sign(array_3_0_io_B_out_sign),
    .io_B_out_exponent(array_3_0_io_B_out_exponent),
    .io_B_out_fraction(array_3_0_io_B_out_fraction),
    .io_C_out_zero(array_3_0_io_C_out_zero),
    .io_C_out_nan(array_3_0_io_C_out_nan),
    .io_C_out_number(array_3_0_io_C_out_number),
    .io_prop_out(array_3_0_io_prop_out)
  );
  logTile array_3_1 ( // @[Array.scala 95:75]
    .clock(array_3_1_clock),
    .io_A_in_zero(array_3_1_io_A_in_zero),
    .io_A_in_nan(array_3_1_io_A_in_nan),
    .io_A_in_sign(array_3_1_io_A_in_sign),
    .io_A_in_exponent(array_3_1_io_A_in_exponent),
    .io_A_in_fraction(array_3_1_io_A_in_fraction),
    .io_B_in_zero(array_3_1_io_B_in_zero),
    .io_B_in_nan(array_3_1_io_B_in_nan),
    .io_B_in_sign(array_3_1_io_B_in_sign),
    .io_B_in_exponent(array_3_1_io_B_in_exponent),
    .io_B_in_fraction(array_3_1_io_B_in_fraction),
    .io_C_in_zero(array_3_1_io_C_in_zero),
    .io_C_in_nan(array_3_1_io_C_in_nan),
    .io_C_in_number(array_3_1_io_C_in_number),
    .io_prop_in(array_3_1_io_prop_in),
    .io_A_out_zero(array_3_1_io_A_out_zero),
    .io_A_out_nan(array_3_1_io_A_out_nan),
    .io_A_out_sign(array_3_1_io_A_out_sign),
    .io_A_out_exponent(array_3_1_io_A_out_exponent),
    .io_A_out_fraction(array_3_1_io_A_out_fraction),
    .io_B_out_zero(array_3_1_io_B_out_zero),
    .io_B_out_nan(array_3_1_io_B_out_nan),
    .io_B_out_sign(array_3_1_io_B_out_sign),
    .io_B_out_exponent(array_3_1_io_B_out_exponent),
    .io_B_out_fraction(array_3_1_io_B_out_fraction),
    .io_C_out_zero(array_3_1_io_C_out_zero),
    .io_C_out_nan(array_3_1_io_C_out_nan),
    .io_C_out_number(array_3_1_io_C_out_number),
    .io_prop_out(array_3_1_io_prop_out)
  );
  logTile array_3_2 ( // @[Array.scala 95:75]
    .clock(array_3_2_clock),
    .io_A_in_zero(array_3_2_io_A_in_zero),
    .io_A_in_nan(array_3_2_io_A_in_nan),
    .io_A_in_sign(array_3_2_io_A_in_sign),
    .io_A_in_exponent(array_3_2_io_A_in_exponent),
    .io_A_in_fraction(array_3_2_io_A_in_fraction),
    .io_B_in_zero(array_3_2_io_B_in_zero),
    .io_B_in_nan(array_3_2_io_B_in_nan),
    .io_B_in_sign(array_3_2_io_B_in_sign),
    .io_B_in_exponent(array_3_2_io_B_in_exponent),
    .io_B_in_fraction(array_3_2_io_B_in_fraction),
    .io_C_in_zero(array_3_2_io_C_in_zero),
    .io_C_in_nan(array_3_2_io_C_in_nan),
    .io_C_in_number(array_3_2_io_C_in_number),
    .io_prop_in(array_3_2_io_prop_in),
    .io_A_out_zero(array_3_2_io_A_out_zero),
    .io_A_out_nan(array_3_2_io_A_out_nan),
    .io_A_out_sign(array_3_2_io_A_out_sign),
    .io_A_out_exponent(array_3_2_io_A_out_exponent),
    .io_A_out_fraction(array_3_2_io_A_out_fraction),
    .io_B_out_zero(array_3_2_io_B_out_zero),
    .io_B_out_nan(array_3_2_io_B_out_nan),
    .io_B_out_sign(array_3_2_io_B_out_sign),
    .io_B_out_exponent(array_3_2_io_B_out_exponent),
    .io_B_out_fraction(array_3_2_io_B_out_fraction),
    .io_C_out_zero(array_3_2_io_C_out_zero),
    .io_C_out_nan(array_3_2_io_C_out_nan),
    .io_C_out_number(array_3_2_io_C_out_number),
    .io_prop_out(array_3_2_io_prop_out)
  );
  logTile array_3_3 ( // @[Array.scala 95:75]
    .clock(array_3_3_clock),
    .io_A_in_zero(array_3_3_io_A_in_zero),
    .io_A_in_nan(array_3_3_io_A_in_nan),
    .io_A_in_sign(array_3_3_io_A_in_sign),
    .io_A_in_exponent(array_3_3_io_A_in_exponent),
    .io_A_in_fraction(array_3_3_io_A_in_fraction),
    .io_B_in_zero(array_3_3_io_B_in_zero),
    .io_B_in_nan(array_3_3_io_B_in_nan),
    .io_B_in_sign(array_3_3_io_B_in_sign),
    .io_B_in_exponent(array_3_3_io_B_in_exponent),
    .io_B_in_fraction(array_3_3_io_B_in_fraction),
    .io_C_in_zero(array_3_3_io_C_in_zero),
    .io_C_in_nan(array_3_3_io_C_in_nan),
    .io_C_in_number(array_3_3_io_C_in_number),
    .io_prop_in(array_3_3_io_prop_in),
    .io_A_out_zero(array_3_3_io_A_out_zero),
    .io_A_out_nan(array_3_3_io_A_out_nan),
    .io_A_out_sign(array_3_3_io_A_out_sign),
    .io_A_out_exponent(array_3_3_io_A_out_exponent),
    .io_A_out_fraction(array_3_3_io_A_out_fraction),
    .io_B_out_zero(array_3_3_io_B_out_zero),
    .io_B_out_nan(array_3_3_io_B_out_nan),
    .io_B_out_sign(array_3_3_io_B_out_sign),
    .io_B_out_exponent(array_3_3_io_B_out_exponent),
    .io_B_out_fraction(array_3_3_io_B_out_fraction),
    .io_C_out_zero(array_3_3_io_C_out_zero),
    .io_C_out_nan(array_3_3_io_C_out_nan),
    .io_C_out_number(array_3_3_io_C_out_number),
    .io_prop_out(array_3_3_io_prop_out)
  );
  toPositUnpacked A_convert_0 ( // @[Array.scala 98:76]
    .io_in(A_convert_0_io_in),
    .io_out_zero(A_convert_0_io_out_zero),
    .io_out_nan(A_convert_0_io_out_nan),
    .io_out_sign(A_convert_0_io_out_sign),
    .io_out_exponent(A_convert_0_io_out_exponent),
    .io_out_fraction(A_convert_0_io_out_fraction)
  );
  toPositUnpacked A_convert_1 ( // @[Array.scala 98:76]
    .io_in(A_convert_1_io_in),
    .io_out_zero(A_convert_1_io_out_zero),
    .io_out_nan(A_convert_1_io_out_nan),
    .io_out_sign(A_convert_1_io_out_sign),
    .io_out_exponent(A_convert_1_io_out_exponent),
    .io_out_fraction(A_convert_1_io_out_fraction)
  );
  toPositUnpacked A_convert_2 ( // @[Array.scala 98:76]
    .io_in(A_convert_2_io_in),
    .io_out_zero(A_convert_2_io_out_zero),
    .io_out_nan(A_convert_2_io_out_nan),
    .io_out_sign(A_convert_2_io_out_sign),
    .io_out_exponent(A_convert_2_io_out_exponent),
    .io_out_fraction(A_convert_2_io_out_fraction)
  );
  toPositUnpacked A_convert_3 ( // @[Array.scala 98:76]
    .io_in(A_convert_3_io_in),
    .io_out_zero(A_convert_3_io_out_zero),
    .io_out_nan(A_convert_3_io_out_nan),
    .io_out_sign(A_convert_3_io_out_sign),
    .io_out_exponent(A_convert_3_io_out_exponent),
    .io_out_fraction(A_convert_3_io_out_fraction)
  );
  toPositUnpacked B_convert_0 ( // @[Array.scala 99:76]
    .io_in(B_convert_0_io_in),
    .io_out_zero(B_convert_0_io_out_zero),
    .io_out_nan(B_convert_0_io_out_nan),
    .io_out_sign(B_convert_0_io_out_sign),
    .io_out_exponent(B_convert_0_io_out_exponent),
    .io_out_fraction(B_convert_0_io_out_fraction)
  );
  toPositUnpacked B_convert_1 ( // @[Array.scala 99:76]
    .io_in(B_convert_1_io_in),
    .io_out_zero(B_convert_1_io_out_zero),
    .io_out_nan(B_convert_1_io_out_nan),
    .io_out_sign(B_convert_1_io_out_sign),
    .io_out_exponent(B_convert_1_io_out_exponent),
    .io_out_fraction(B_convert_1_io_out_fraction)
  );
  toPositUnpacked B_convert_2 ( // @[Array.scala 99:76]
    .io_in(B_convert_2_io_in),
    .io_out_zero(B_convert_2_io_out_zero),
    .io_out_nan(B_convert_2_io_out_nan),
    .io_out_sign(B_convert_2_io_out_sign),
    .io_out_exponent(B_convert_2_io_out_exponent),
    .io_out_fraction(B_convert_2_io_out_fraction)
  );
  toPositUnpacked B_convert_3 ( // @[Array.scala 99:76]
    .io_in(B_convert_3_io_in),
    .io_out_zero(B_convert_3_io_out_zero),
    .io_out_nan(B_convert_3_io_out_nan),
    .io_out_sign(B_convert_3_io_out_sign),
    .io_out_exponent(B_convert_3_io_out_exponent),
    .io_out_fraction(B_convert_3_io_out_fraction)
  );
  assign io_C_out_0_zero = array_3_0_io_C_out_zero; // @[Array.scala 111:37]
  assign io_C_out_0_nan = array_3_0_io_C_out_nan; // @[Array.scala 111:37]
  assign io_C_out_0_number = array_3_0_io_C_out_number; // @[Array.scala 111:37]
  assign io_C_out_1_zero = array_3_1_io_C_out_zero; // @[Array.scala 111:37]
  assign io_C_out_1_nan = array_3_1_io_C_out_nan; // @[Array.scala 111:37]
  assign io_C_out_1_number = array_3_1_io_C_out_number; // @[Array.scala 111:37]
  assign io_C_out_2_zero = array_3_2_io_C_out_zero; // @[Array.scala 111:37]
  assign io_C_out_2_nan = array_3_2_io_C_out_nan; // @[Array.scala 111:37]
  assign io_C_out_2_number = array_3_2_io_C_out_number; // @[Array.scala 111:37]
  assign io_C_out_3_zero = array_3_3_io_C_out_zero; // @[Array.scala 111:37]
  assign io_C_out_3_nan = array_3_3_io_C_out_nan; // @[Array.scala 111:37]
  assign io_C_out_3_number = array_3_3_io_C_out_number; // @[Array.scala 111:37]
  assign array_0_0_clock = clock;
  assign array_0_0_io_A_in_zero = A_convert_0_io_out_zero; // @[Array.scala 103:45]
  assign array_0_0_io_A_in_nan = A_convert_0_io_out_nan; // @[Array.scala 103:45]
  assign array_0_0_io_A_in_sign = A_convert_0_io_out_sign; // @[Array.scala 103:45]
  assign array_0_0_io_A_in_exponent = A_convert_0_io_out_exponent; // @[Array.scala 103:45]
  assign array_0_0_io_A_in_fraction = A_convert_0_io_out_fraction; // @[Array.scala 103:45]
  assign array_0_0_io_B_in_zero = B_convert_0_io_out_zero; // @[Array.scala 116:45]
  assign array_0_0_io_B_in_nan = B_convert_0_io_out_nan; // @[Array.scala 116:45]
  assign array_0_0_io_B_in_sign = B_convert_0_io_out_sign; // @[Array.scala 116:45]
  assign array_0_0_io_B_in_exponent = B_convert_0_io_out_exponent; // @[Array.scala 116:45]
  assign array_0_0_io_B_in_fraction = B_convert_0_io_out_fraction; // @[Array.scala 116:45]
  assign array_0_0_io_C_in_zero = io_C_in_0_zero; // @[Array.scala 104:45]
  assign array_0_0_io_C_in_nan = io_C_in_0_nan; // @[Array.scala 104:45]
  assign array_0_0_io_C_in_number = io_C_in_0_number; // @[Array.scala 104:45]
  assign array_0_0_io_prop_in = io_prop_in_0; // @[Array.scala 105:48]
  assign array_0_1_clock = clock;
  assign array_0_1_io_A_in_zero = A_convert_1_io_out_zero; // @[Array.scala 103:45]
  assign array_0_1_io_A_in_nan = A_convert_1_io_out_nan; // @[Array.scala 103:45]
  assign array_0_1_io_A_in_sign = A_convert_1_io_out_sign; // @[Array.scala 103:45]
  assign array_0_1_io_A_in_exponent = A_convert_1_io_out_exponent; // @[Array.scala 103:45]
  assign array_0_1_io_A_in_fraction = A_convert_1_io_out_fraction; // @[Array.scala 103:45]
  assign array_0_1_io_B_in_zero = array_0_0_io_B_out_zero; // @[Array.scala 118:53]
  assign array_0_1_io_B_in_nan = array_0_0_io_B_out_nan; // @[Array.scala 118:53]
  assign array_0_1_io_B_in_sign = array_0_0_io_B_out_sign; // @[Array.scala 118:53]
  assign array_0_1_io_B_in_exponent = array_0_0_io_B_out_exponent; // @[Array.scala 118:53]
  assign array_0_1_io_B_in_fraction = array_0_0_io_B_out_fraction; // @[Array.scala 118:53]
  assign array_0_1_io_C_in_zero = io_C_in_1_zero; // @[Array.scala 104:45]
  assign array_0_1_io_C_in_nan = io_C_in_1_nan; // @[Array.scala 104:45]
  assign array_0_1_io_C_in_number = io_C_in_1_number; // @[Array.scala 104:45]
  assign array_0_1_io_prop_in = io_prop_in_1; // @[Array.scala 105:48]
  assign array_0_2_clock = clock;
  assign array_0_2_io_A_in_zero = A_convert_2_io_out_zero; // @[Array.scala 103:45]
  assign array_0_2_io_A_in_nan = A_convert_2_io_out_nan; // @[Array.scala 103:45]
  assign array_0_2_io_A_in_sign = A_convert_2_io_out_sign; // @[Array.scala 103:45]
  assign array_0_2_io_A_in_exponent = A_convert_2_io_out_exponent; // @[Array.scala 103:45]
  assign array_0_2_io_A_in_fraction = A_convert_2_io_out_fraction; // @[Array.scala 103:45]
  assign array_0_2_io_B_in_zero = array_0_1_io_B_out_zero; // @[Array.scala 118:53]
  assign array_0_2_io_B_in_nan = array_0_1_io_B_out_nan; // @[Array.scala 118:53]
  assign array_0_2_io_B_in_sign = array_0_1_io_B_out_sign; // @[Array.scala 118:53]
  assign array_0_2_io_B_in_exponent = array_0_1_io_B_out_exponent; // @[Array.scala 118:53]
  assign array_0_2_io_B_in_fraction = array_0_1_io_B_out_fraction; // @[Array.scala 118:53]
  assign array_0_2_io_C_in_zero = io_C_in_2_zero; // @[Array.scala 104:45]
  assign array_0_2_io_C_in_nan = io_C_in_2_nan; // @[Array.scala 104:45]
  assign array_0_2_io_C_in_number = io_C_in_2_number; // @[Array.scala 104:45]
  assign array_0_2_io_prop_in = io_prop_in_2; // @[Array.scala 105:48]
  assign array_0_3_clock = clock;
  assign array_0_3_io_A_in_zero = A_convert_3_io_out_zero; // @[Array.scala 103:45]
  assign array_0_3_io_A_in_nan = A_convert_3_io_out_nan; // @[Array.scala 103:45]
  assign array_0_3_io_A_in_sign = A_convert_3_io_out_sign; // @[Array.scala 103:45]
  assign array_0_3_io_A_in_exponent = A_convert_3_io_out_exponent; // @[Array.scala 103:45]
  assign array_0_3_io_A_in_fraction = A_convert_3_io_out_fraction; // @[Array.scala 103:45]
  assign array_0_3_io_B_in_zero = array_0_2_io_B_out_zero; // @[Array.scala 118:53]
  assign array_0_3_io_B_in_nan = array_0_2_io_B_out_nan; // @[Array.scala 118:53]
  assign array_0_3_io_B_in_sign = array_0_2_io_B_out_sign; // @[Array.scala 118:53]
  assign array_0_3_io_B_in_exponent = array_0_2_io_B_out_exponent; // @[Array.scala 118:53]
  assign array_0_3_io_B_in_fraction = array_0_2_io_B_out_fraction; // @[Array.scala 118:53]
  assign array_0_3_io_C_in_zero = io_C_in_3_zero; // @[Array.scala 104:45]
  assign array_0_3_io_C_in_nan = io_C_in_3_nan; // @[Array.scala 104:45]
  assign array_0_3_io_C_in_number = io_C_in_3_number; // @[Array.scala 104:45]
  assign array_0_3_io_prop_in = io_prop_in_3; // @[Array.scala 105:48]
  assign array_1_0_clock = clock;
  assign array_1_0_io_A_in_zero = array_0_0_io_A_out_zero; // @[Array.scala 107:53]
  assign array_1_0_io_A_in_nan = array_0_0_io_A_out_nan; // @[Array.scala 107:53]
  assign array_1_0_io_A_in_sign = array_0_0_io_A_out_sign; // @[Array.scala 107:53]
  assign array_1_0_io_A_in_exponent = array_0_0_io_A_out_exponent; // @[Array.scala 107:53]
  assign array_1_0_io_A_in_fraction = array_0_0_io_A_out_fraction; // @[Array.scala 107:53]
  assign array_1_0_io_B_in_zero = B_convert_1_io_out_zero; // @[Array.scala 116:45]
  assign array_1_0_io_B_in_nan = B_convert_1_io_out_nan; // @[Array.scala 116:45]
  assign array_1_0_io_B_in_sign = B_convert_1_io_out_sign; // @[Array.scala 116:45]
  assign array_1_0_io_B_in_exponent = B_convert_1_io_out_exponent; // @[Array.scala 116:45]
  assign array_1_0_io_B_in_fraction = B_convert_1_io_out_fraction; // @[Array.scala 116:45]
  assign array_1_0_io_C_in_zero = array_0_0_io_C_out_zero; // @[Array.scala 108:53]
  assign array_1_0_io_C_in_nan = array_0_0_io_C_out_nan; // @[Array.scala 108:53]
  assign array_1_0_io_C_in_number = array_0_0_io_C_out_number; // @[Array.scala 108:53]
  assign array_1_0_io_prop_in = array_0_0_io_prop_out; // @[Array.scala 109:56]
  assign array_1_1_clock = clock;
  assign array_1_1_io_A_in_zero = array_0_1_io_A_out_zero; // @[Array.scala 107:53]
  assign array_1_1_io_A_in_nan = array_0_1_io_A_out_nan; // @[Array.scala 107:53]
  assign array_1_1_io_A_in_sign = array_0_1_io_A_out_sign; // @[Array.scala 107:53]
  assign array_1_1_io_A_in_exponent = array_0_1_io_A_out_exponent; // @[Array.scala 107:53]
  assign array_1_1_io_A_in_fraction = array_0_1_io_A_out_fraction; // @[Array.scala 107:53]
  assign array_1_1_io_B_in_zero = array_1_0_io_B_out_zero; // @[Array.scala 118:53]
  assign array_1_1_io_B_in_nan = array_1_0_io_B_out_nan; // @[Array.scala 118:53]
  assign array_1_1_io_B_in_sign = array_1_0_io_B_out_sign; // @[Array.scala 118:53]
  assign array_1_1_io_B_in_exponent = array_1_0_io_B_out_exponent; // @[Array.scala 118:53]
  assign array_1_1_io_B_in_fraction = array_1_0_io_B_out_fraction; // @[Array.scala 118:53]
  assign array_1_1_io_C_in_zero = array_0_1_io_C_out_zero; // @[Array.scala 108:53]
  assign array_1_1_io_C_in_nan = array_0_1_io_C_out_nan; // @[Array.scala 108:53]
  assign array_1_1_io_C_in_number = array_0_1_io_C_out_number; // @[Array.scala 108:53]
  assign array_1_1_io_prop_in = array_0_1_io_prop_out; // @[Array.scala 109:56]
  assign array_1_2_clock = clock;
  assign array_1_2_io_A_in_zero = array_0_2_io_A_out_zero; // @[Array.scala 107:53]
  assign array_1_2_io_A_in_nan = array_0_2_io_A_out_nan; // @[Array.scala 107:53]
  assign array_1_2_io_A_in_sign = array_0_2_io_A_out_sign; // @[Array.scala 107:53]
  assign array_1_2_io_A_in_exponent = array_0_2_io_A_out_exponent; // @[Array.scala 107:53]
  assign array_1_2_io_A_in_fraction = array_0_2_io_A_out_fraction; // @[Array.scala 107:53]
  assign array_1_2_io_B_in_zero = array_1_1_io_B_out_zero; // @[Array.scala 118:53]
  assign array_1_2_io_B_in_nan = array_1_1_io_B_out_nan; // @[Array.scala 118:53]
  assign array_1_2_io_B_in_sign = array_1_1_io_B_out_sign; // @[Array.scala 118:53]
  assign array_1_2_io_B_in_exponent = array_1_1_io_B_out_exponent; // @[Array.scala 118:53]
  assign array_1_2_io_B_in_fraction = array_1_1_io_B_out_fraction; // @[Array.scala 118:53]
  assign array_1_2_io_C_in_zero = array_0_2_io_C_out_zero; // @[Array.scala 108:53]
  assign array_1_2_io_C_in_nan = array_0_2_io_C_out_nan; // @[Array.scala 108:53]
  assign array_1_2_io_C_in_number = array_0_2_io_C_out_number; // @[Array.scala 108:53]
  assign array_1_2_io_prop_in = array_0_2_io_prop_out; // @[Array.scala 109:56]
  assign array_1_3_clock = clock;
  assign array_1_3_io_A_in_zero = array_0_3_io_A_out_zero; // @[Array.scala 107:53]
  assign array_1_3_io_A_in_nan = array_0_3_io_A_out_nan; // @[Array.scala 107:53]
  assign array_1_3_io_A_in_sign = array_0_3_io_A_out_sign; // @[Array.scala 107:53]
  assign array_1_3_io_A_in_exponent = array_0_3_io_A_out_exponent; // @[Array.scala 107:53]
  assign array_1_3_io_A_in_fraction = array_0_3_io_A_out_fraction; // @[Array.scala 107:53]
  assign array_1_3_io_B_in_zero = array_1_2_io_B_out_zero; // @[Array.scala 118:53]
  assign array_1_3_io_B_in_nan = array_1_2_io_B_out_nan; // @[Array.scala 118:53]
  assign array_1_3_io_B_in_sign = array_1_2_io_B_out_sign; // @[Array.scala 118:53]
  assign array_1_3_io_B_in_exponent = array_1_2_io_B_out_exponent; // @[Array.scala 118:53]
  assign array_1_3_io_B_in_fraction = array_1_2_io_B_out_fraction; // @[Array.scala 118:53]
  assign array_1_3_io_C_in_zero = array_0_3_io_C_out_zero; // @[Array.scala 108:53]
  assign array_1_3_io_C_in_nan = array_0_3_io_C_out_nan; // @[Array.scala 108:53]
  assign array_1_3_io_C_in_number = array_0_3_io_C_out_number; // @[Array.scala 108:53]
  assign array_1_3_io_prop_in = array_0_3_io_prop_out; // @[Array.scala 109:56]
  assign array_2_0_clock = clock;
  assign array_2_0_io_A_in_zero = array_1_0_io_A_out_zero; // @[Array.scala 107:53]
  assign array_2_0_io_A_in_nan = array_1_0_io_A_out_nan; // @[Array.scala 107:53]
  assign array_2_0_io_A_in_sign = array_1_0_io_A_out_sign; // @[Array.scala 107:53]
  assign array_2_0_io_A_in_exponent = array_1_0_io_A_out_exponent; // @[Array.scala 107:53]
  assign array_2_0_io_A_in_fraction = array_1_0_io_A_out_fraction; // @[Array.scala 107:53]
  assign array_2_0_io_B_in_zero = B_convert_2_io_out_zero; // @[Array.scala 116:45]
  assign array_2_0_io_B_in_nan = B_convert_2_io_out_nan; // @[Array.scala 116:45]
  assign array_2_0_io_B_in_sign = B_convert_2_io_out_sign; // @[Array.scala 116:45]
  assign array_2_0_io_B_in_exponent = B_convert_2_io_out_exponent; // @[Array.scala 116:45]
  assign array_2_0_io_B_in_fraction = B_convert_2_io_out_fraction; // @[Array.scala 116:45]
  assign array_2_0_io_C_in_zero = array_1_0_io_C_out_zero; // @[Array.scala 108:53]
  assign array_2_0_io_C_in_nan = array_1_0_io_C_out_nan; // @[Array.scala 108:53]
  assign array_2_0_io_C_in_number = array_1_0_io_C_out_number; // @[Array.scala 108:53]
  assign array_2_0_io_prop_in = array_1_0_io_prop_out; // @[Array.scala 109:56]
  assign array_2_1_clock = clock;
  assign array_2_1_io_A_in_zero = array_1_1_io_A_out_zero; // @[Array.scala 107:53]
  assign array_2_1_io_A_in_nan = array_1_1_io_A_out_nan; // @[Array.scala 107:53]
  assign array_2_1_io_A_in_sign = array_1_1_io_A_out_sign; // @[Array.scala 107:53]
  assign array_2_1_io_A_in_exponent = array_1_1_io_A_out_exponent; // @[Array.scala 107:53]
  assign array_2_1_io_A_in_fraction = array_1_1_io_A_out_fraction; // @[Array.scala 107:53]
  assign array_2_1_io_B_in_zero = array_2_0_io_B_out_zero; // @[Array.scala 118:53]
  assign array_2_1_io_B_in_nan = array_2_0_io_B_out_nan; // @[Array.scala 118:53]
  assign array_2_1_io_B_in_sign = array_2_0_io_B_out_sign; // @[Array.scala 118:53]
  assign array_2_1_io_B_in_exponent = array_2_0_io_B_out_exponent; // @[Array.scala 118:53]
  assign array_2_1_io_B_in_fraction = array_2_0_io_B_out_fraction; // @[Array.scala 118:53]
  assign array_2_1_io_C_in_zero = array_1_1_io_C_out_zero; // @[Array.scala 108:53]
  assign array_2_1_io_C_in_nan = array_1_1_io_C_out_nan; // @[Array.scala 108:53]
  assign array_2_1_io_C_in_number = array_1_1_io_C_out_number; // @[Array.scala 108:53]
  assign array_2_1_io_prop_in = array_1_1_io_prop_out; // @[Array.scala 109:56]
  assign array_2_2_clock = clock;
  assign array_2_2_io_A_in_zero = array_1_2_io_A_out_zero; // @[Array.scala 107:53]
  assign array_2_2_io_A_in_nan = array_1_2_io_A_out_nan; // @[Array.scala 107:53]
  assign array_2_2_io_A_in_sign = array_1_2_io_A_out_sign; // @[Array.scala 107:53]
  assign array_2_2_io_A_in_exponent = array_1_2_io_A_out_exponent; // @[Array.scala 107:53]
  assign array_2_2_io_A_in_fraction = array_1_2_io_A_out_fraction; // @[Array.scala 107:53]
  assign array_2_2_io_B_in_zero = array_2_1_io_B_out_zero; // @[Array.scala 118:53]
  assign array_2_2_io_B_in_nan = array_2_1_io_B_out_nan; // @[Array.scala 118:53]
  assign array_2_2_io_B_in_sign = array_2_1_io_B_out_sign; // @[Array.scala 118:53]
  assign array_2_2_io_B_in_exponent = array_2_1_io_B_out_exponent; // @[Array.scala 118:53]
  assign array_2_2_io_B_in_fraction = array_2_1_io_B_out_fraction; // @[Array.scala 118:53]
  assign array_2_2_io_C_in_zero = array_1_2_io_C_out_zero; // @[Array.scala 108:53]
  assign array_2_2_io_C_in_nan = array_1_2_io_C_out_nan; // @[Array.scala 108:53]
  assign array_2_2_io_C_in_number = array_1_2_io_C_out_number; // @[Array.scala 108:53]
  assign array_2_2_io_prop_in = array_1_2_io_prop_out; // @[Array.scala 109:56]
  assign array_2_3_clock = clock;
  assign array_2_3_io_A_in_zero = array_1_3_io_A_out_zero; // @[Array.scala 107:53]
  assign array_2_3_io_A_in_nan = array_1_3_io_A_out_nan; // @[Array.scala 107:53]
  assign array_2_3_io_A_in_sign = array_1_3_io_A_out_sign; // @[Array.scala 107:53]
  assign array_2_3_io_A_in_exponent = array_1_3_io_A_out_exponent; // @[Array.scala 107:53]
  assign array_2_3_io_A_in_fraction = array_1_3_io_A_out_fraction; // @[Array.scala 107:53]
  assign array_2_3_io_B_in_zero = array_2_2_io_B_out_zero; // @[Array.scala 118:53]
  assign array_2_3_io_B_in_nan = array_2_2_io_B_out_nan; // @[Array.scala 118:53]
  assign array_2_3_io_B_in_sign = array_2_2_io_B_out_sign; // @[Array.scala 118:53]
  assign array_2_3_io_B_in_exponent = array_2_2_io_B_out_exponent; // @[Array.scala 118:53]
  assign array_2_3_io_B_in_fraction = array_2_2_io_B_out_fraction; // @[Array.scala 118:53]
  assign array_2_3_io_C_in_zero = array_1_3_io_C_out_zero; // @[Array.scala 108:53]
  assign array_2_3_io_C_in_nan = array_1_3_io_C_out_nan; // @[Array.scala 108:53]
  assign array_2_3_io_C_in_number = array_1_3_io_C_out_number; // @[Array.scala 108:53]
  assign array_2_3_io_prop_in = array_1_3_io_prop_out; // @[Array.scala 109:56]
  assign array_3_0_clock = clock;
  assign array_3_0_io_A_in_zero = array_2_0_io_A_out_zero; // @[Array.scala 107:53]
  assign array_3_0_io_A_in_nan = array_2_0_io_A_out_nan; // @[Array.scala 107:53]
  assign array_3_0_io_A_in_sign = array_2_0_io_A_out_sign; // @[Array.scala 107:53]
  assign array_3_0_io_A_in_exponent = array_2_0_io_A_out_exponent; // @[Array.scala 107:53]
  assign array_3_0_io_A_in_fraction = array_2_0_io_A_out_fraction; // @[Array.scala 107:53]
  assign array_3_0_io_B_in_zero = B_convert_3_io_out_zero; // @[Array.scala 116:45]
  assign array_3_0_io_B_in_nan = B_convert_3_io_out_nan; // @[Array.scala 116:45]
  assign array_3_0_io_B_in_sign = B_convert_3_io_out_sign; // @[Array.scala 116:45]
  assign array_3_0_io_B_in_exponent = B_convert_3_io_out_exponent; // @[Array.scala 116:45]
  assign array_3_0_io_B_in_fraction = B_convert_3_io_out_fraction; // @[Array.scala 116:45]
  assign array_3_0_io_C_in_zero = array_2_0_io_C_out_zero; // @[Array.scala 108:53]
  assign array_3_0_io_C_in_nan = array_2_0_io_C_out_nan; // @[Array.scala 108:53]
  assign array_3_0_io_C_in_number = array_2_0_io_C_out_number; // @[Array.scala 108:53]
  assign array_3_0_io_prop_in = array_2_0_io_prop_out; // @[Array.scala 109:56]
  assign array_3_1_clock = clock;
  assign array_3_1_io_A_in_zero = array_2_1_io_A_out_zero; // @[Array.scala 107:53]
  assign array_3_1_io_A_in_nan = array_2_1_io_A_out_nan; // @[Array.scala 107:53]
  assign array_3_1_io_A_in_sign = array_2_1_io_A_out_sign; // @[Array.scala 107:53]
  assign array_3_1_io_A_in_exponent = array_2_1_io_A_out_exponent; // @[Array.scala 107:53]
  assign array_3_1_io_A_in_fraction = array_2_1_io_A_out_fraction; // @[Array.scala 107:53]
  assign array_3_1_io_B_in_zero = array_3_0_io_B_out_zero; // @[Array.scala 118:53]
  assign array_3_1_io_B_in_nan = array_3_0_io_B_out_nan; // @[Array.scala 118:53]
  assign array_3_1_io_B_in_sign = array_3_0_io_B_out_sign; // @[Array.scala 118:53]
  assign array_3_1_io_B_in_exponent = array_3_0_io_B_out_exponent; // @[Array.scala 118:53]
  assign array_3_1_io_B_in_fraction = array_3_0_io_B_out_fraction; // @[Array.scala 118:53]
  assign array_3_1_io_C_in_zero = array_2_1_io_C_out_zero; // @[Array.scala 108:53]
  assign array_3_1_io_C_in_nan = array_2_1_io_C_out_nan; // @[Array.scala 108:53]
  assign array_3_1_io_C_in_number = array_2_1_io_C_out_number; // @[Array.scala 108:53]
  assign array_3_1_io_prop_in = array_2_1_io_prop_out; // @[Array.scala 109:56]
  assign array_3_2_clock = clock;
  assign array_3_2_io_A_in_zero = array_2_2_io_A_out_zero; // @[Array.scala 107:53]
  assign array_3_2_io_A_in_nan = array_2_2_io_A_out_nan; // @[Array.scala 107:53]
  assign array_3_2_io_A_in_sign = array_2_2_io_A_out_sign; // @[Array.scala 107:53]
  assign array_3_2_io_A_in_exponent = array_2_2_io_A_out_exponent; // @[Array.scala 107:53]
  assign array_3_2_io_A_in_fraction = array_2_2_io_A_out_fraction; // @[Array.scala 107:53]
  assign array_3_2_io_B_in_zero = array_3_1_io_B_out_zero; // @[Array.scala 118:53]
  assign array_3_2_io_B_in_nan = array_3_1_io_B_out_nan; // @[Array.scala 118:53]
  assign array_3_2_io_B_in_sign = array_3_1_io_B_out_sign; // @[Array.scala 118:53]
  assign array_3_2_io_B_in_exponent = array_3_1_io_B_out_exponent; // @[Array.scala 118:53]
  assign array_3_2_io_B_in_fraction = array_3_1_io_B_out_fraction; // @[Array.scala 118:53]
  assign array_3_2_io_C_in_zero = array_2_2_io_C_out_zero; // @[Array.scala 108:53]
  assign array_3_2_io_C_in_nan = array_2_2_io_C_out_nan; // @[Array.scala 108:53]
  assign array_3_2_io_C_in_number = array_2_2_io_C_out_number; // @[Array.scala 108:53]
  assign array_3_2_io_prop_in = array_2_2_io_prop_out; // @[Array.scala 109:56]
  assign array_3_3_clock = clock;
  assign array_3_3_io_A_in_zero = array_2_3_io_A_out_zero; // @[Array.scala 107:53]
  assign array_3_3_io_A_in_nan = array_2_3_io_A_out_nan; // @[Array.scala 107:53]
  assign array_3_3_io_A_in_sign = array_2_3_io_A_out_sign; // @[Array.scala 107:53]
  assign array_3_3_io_A_in_exponent = array_2_3_io_A_out_exponent; // @[Array.scala 107:53]
  assign array_3_3_io_A_in_fraction = array_2_3_io_A_out_fraction; // @[Array.scala 107:53]
  assign array_3_3_io_B_in_zero = array_3_2_io_B_out_zero; // @[Array.scala 118:53]
  assign array_3_3_io_B_in_nan = array_3_2_io_B_out_nan; // @[Array.scala 118:53]
  assign array_3_3_io_B_in_sign = array_3_2_io_B_out_sign; // @[Array.scala 118:53]
  assign array_3_3_io_B_in_exponent = array_3_2_io_B_out_exponent; // @[Array.scala 118:53]
  assign array_3_3_io_B_in_fraction = array_3_2_io_B_out_fraction; // @[Array.scala 118:53]
  assign array_3_3_io_C_in_zero = array_2_3_io_C_out_zero; // @[Array.scala 108:53]
  assign array_3_3_io_C_in_nan = array_2_3_io_C_out_nan; // @[Array.scala 108:53]
  assign array_3_3_io_C_in_number = array_2_3_io_C_out_number; // @[Array.scala 108:53]
  assign array_3_3_io_prop_in = array_2_3_io_prop_out; // @[Array.scala 109:56]
  assign A_convert_0_io_in = io_A_in_0; // @[Array.scala 102:44]
  assign A_convert_1_io_in = io_A_in_1; // @[Array.scala 102:44]
  assign A_convert_2_io_in = io_A_in_2; // @[Array.scala 102:44]
  assign A_convert_3_io_in = io_A_in_3; // @[Array.scala 102:44]
  assign B_convert_0_io_in = io_B_in_0; // @[Array.scala 115:44]
  assign B_convert_1_io_in = io_B_in_1; // @[Array.scala 115:44]
  assign B_convert_2_io_in = io_B_in_2; // @[Array.scala 115:44]
  assign B_convert_3_io_in = io_B_in_3; // @[Array.scala 115:44]
endmodule
