module toPositUnpacked(
  input         clock,
  input         reset,
  input  [15:0] io_in,
  output        io_out_sign,
  output [27:0] io_out_exponent,
  output [11:0] io_out_fraction
);
  wire [14:0] _T_3; // @[Bitwise.scala 71:12]
  wire [14:0] _T_4; // @[Conversion.scala 16:48]
  wire [14:0] _GEN_0; // @[Conversion.scala 16:85]
  wire [14:0] others; // @[Conversion.scala 16:85]
  wire [14:0] _T_7; // @[Conversion.scala 17:122]
  wire [7:0] _T_12; // @[Bitwise.scala 102:31]
  wire [7:0] _T_14; // @[Bitwise.scala 102:65]
  wire [7:0] _T_16; // @[Bitwise.scala 102:75]
  wire [7:0] _T_17; // @[Bitwise.scala 102:39]
  wire [7:0] _GEN_1; // @[Bitwise.scala 102:31]
  wire [7:0] _T_22; // @[Bitwise.scala 102:31]
  wire [7:0] _T_24; // @[Bitwise.scala 102:65]
  wire [7:0] _T_26; // @[Bitwise.scala 102:75]
  wire [7:0] _T_27; // @[Bitwise.scala 102:39]
  wire [7:0] _GEN_2; // @[Bitwise.scala 102:31]
  wire [7:0] _T_32; // @[Bitwise.scala 102:31]
  wire [7:0] _T_34; // @[Bitwise.scala 102:65]
  wire [7:0] _T_36; // @[Bitwise.scala 102:75]
  wire [7:0] _T_37; // @[Bitwise.scala 102:39]
  wire [14:0] _T_57; // @[Cat.scala 29:58]
  wire [3:0] _T_73; // @[Mux.scala 47:69]
  wire [3:0] _T_74; // @[Mux.scala 47:69]
  wire [3:0] _T_75; // @[Mux.scala 47:69]
  wire [3:0] _T_76; // @[Mux.scala 47:69]
  wire [3:0] _T_77; // @[Mux.scala 47:69]
  wire [3:0] _T_78; // @[Mux.scala 47:69]
  wire [3:0] _T_79; // @[Mux.scala 47:69]
  wire [3:0] _T_80; // @[Mux.scala 47:69]
  wire [3:0] _T_81; // @[Mux.scala 47:69]
  wire [3:0] _T_82; // @[Mux.scala 47:69]
  wire [3:0] _T_83; // @[Mux.scala 47:69]
  wire [3:0] _T_84; // @[Mux.scala 47:69]
  wire [3:0] _T_85; // @[Mux.scala 47:69]
  wire [3:0] regime; // @[Mux.scala 47:69]
  assign _T_3 = io_out_sign ? 15'h7fff : 15'h0; // @[Bitwise.scala 71:12]
  assign _T_4 = io_in[14:0] ^ _T_3; // @[Conversion.scala 16:48]
  assign _GEN_0 = {{14'd0}, io_out_sign}; // @[Conversion.scala 16:85]
  assign others = _T_4 + _GEN_0; // @[Conversion.scala 16:85]
  assign _T_7 = ~others; // @[Conversion.scala 17:122]
  assign _T_12 = {{4'd0}, _T_7[7:4]}; // @[Bitwise.scala 102:31]
  assign _T_14 = {_T_7[3:0], 4'h0}; // @[Bitwise.scala 102:65]
  assign _T_16 = _T_14 & 8'hf0; // @[Bitwise.scala 102:75]
  assign _T_17 = _T_12 | _T_16; // @[Bitwise.scala 102:39]
  assign _GEN_1 = {{2'd0}, _T_17[7:2]}; // @[Bitwise.scala 102:31]
  assign _T_22 = _GEN_1 & 8'h33; // @[Bitwise.scala 102:31]
  assign _T_24 = {_T_17[5:0], 2'h0}; // @[Bitwise.scala 102:65]
  assign _T_26 = _T_24 & 8'hcc; // @[Bitwise.scala 102:75]
  assign _T_27 = _T_22 | _T_26; // @[Bitwise.scala 102:39]
  assign _GEN_2 = {{1'd0}, _T_27[7:1]}; // @[Bitwise.scala 102:31]
  assign _T_32 = _GEN_2 & 8'h55; // @[Bitwise.scala 102:31]
  assign _T_34 = {_T_27[6:0], 1'h0}; // @[Bitwise.scala 102:65]
  assign _T_36 = _T_34 & 8'haa; // @[Bitwise.scala 102:75]
  assign _T_37 = _T_32 | _T_36; // @[Bitwise.scala 102:39]
  assign _T_57 = {_T_37,_T_7[8],_T_7[9],_T_7[10],_T_7[11],_T_7[12],_T_7[13],_T_7[14]}; // @[Cat.scala 29:58]
  assign _T_73 = _T_57[13] ? 4'hd : 4'he; // @[Mux.scala 47:69]
  assign _T_74 = _T_57[12] ? 4'hc : _T_73; // @[Mux.scala 47:69]
  assign _T_75 = _T_57[11] ? 4'hb : _T_74; // @[Mux.scala 47:69]
  assign _T_76 = _T_57[10] ? 4'ha : _T_75; // @[Mux.scala 47:69]
  assign _T_77 = _T_57[9] ? 4'h9 : _T_76; // @[Mux.scala 47:69]
  assign _T_78 = _T_57[8] ? 4'h8 : _T_77; // @[Mux.scala 47:69]
  assign _T_79 = _T_57[7] ? 4'h7 : _T_78; // @[Mux.scala 47:69]
  assign _T_80 = _T_57[6] ? 4'h6 : _T_79; // @[Mux.scala 47:69]
  assign _T_81 = _T_57[5] ? 4'h5 : _T_80; // @[Mux.scala 47:69]
  assign _T_82 = _T_57[4] ? 4'h4 : _T_81; // @[Mux.scala 47:69]
  assign _T_83 = _T_57[3] ? 4'h3 : _T_82; // @[Mux.scala 47:69]
  assign _T_84 = _T_57[2] ? 4'h2 : _T_83; // @[Mux.scala 47:69]
  assign _T_85 = _T_57[1] ? 4'h1 : _T_84; // @[Mux.scala 47:69]
  assign regime = _T_57[0] ? 4'h0 : _T_85; // @[Mux.scala 47:69]
  assign io_out_sign = io_in[15]; // @[Conversion.scala 14:21]
  assign io_out_exponent = {{24'd0}, regime}; // @[Conversion.scala 18:25]
  assign io_out_fraction = 12'h0; // @[Conversion.scala 19:25]
endmodule
